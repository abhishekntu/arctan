--------------------------------------------------------------------------------
--                             LZOC_14_F400_uid4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOC_14_F400_uid4 is
   port ( clk, rst : in std_logic;
          I : in  std_logic_vector(13 downto 0);
          OZB : in  std_logic;
          O : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of LZOC_14_F400_uid4 is
signal sozb, sozb_d1, sozb_d2 :  std_logic;
signal level4 :  std_logic_vector(15 downto 0);
signal digit4, digit4_d1, digit4_d2 :  std_logic;
signal level3, level3_d1 :  std_logic_vector(7 downto 0);
signal digit3, digit3_d1 :  std_logic;
signal level2 :  std_logic_vector(3 downto 0);
signal digit2, digit2_d1 :  std_logic;
signal level1, level1_d1 :  std_logic_vector(1 downto 0);
signal digit1 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sozb_d1 <=  sozb;
            sozb_d2 <=  sozb_d1;
            digit4_d1 <=  digit4;
            digit4_d2 <=  digit4_d1;
            level3_d1 <=  level3;
            digit3_d1 <=  digit3;
            digit2_d1 <=  digit2;
            level1_d1 <=  level1;
         end if;
      end process;
   sozb <= OZB;
   level4<= I& (1 downto 0 => not(sozb));
   digit4<= '1' when level4(15 downto 8) = (15 downto 8 => sozb) else '0';
   level3<= level4(7 downto 0) when digit4='1' else level4(15 downto 8);
   ----------------Synchro barrier, entering cycle 1----------------
   digit3<= '1' when level3_d1(7 downto 4) = (7 downto 4 => sozb_d1) else '0';
   level2<= level3_d1(3 downto 0) when digit3='1' else level3_d1(7 downto 4);
   digit2<= '1' when level2(3 downto 2) = (3 downto 2 => sozb_d1) else '0';
   level1<= level2(1 downto 0) when digit2='1' else level2(3 downto 2);
   ----------------Synchro barrier, entering cycle 2----------------
   digit1<= '1' when level1_d1(1 downto 1) = (1 downto 1 => sozb_d2) else '0';
   O <= digit4_d2 & digit3_d1 & digit2_d1 & digit1;
end architecture;

--------------------------------------------------------------------------------
--                     LeftShifter_15_by_max_14_F400_uid8
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter_15_by_max_14_F400_uid8 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(14 downto 0);
          S : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(28 downto 0)   );
end entity;

architecture arch of LeftShifter_15_by_max_14_F400_uid8 is
signal level0 :  std_logic_vector(14 downto 0);
signal ps, ps_d1 :  std_logic_vector(3 downto 0);
signal level1 :  std_logic_vector(15 downto 0);
signal level2 :  std_logic_vector(17 downto 0);
signal level3, level3_d1 :  std_logic_vector(21 downto 0);
signal level4 :  std_logic_vector(29 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            level3_d1 <=  level3;
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<= level0 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => '0') & level0;
   level2<= level1 & (1 downto 0 => '0') when ps(1)= '1' else     (1 downto 0 => '0') & level1;
   level3<= level2 & (3 downto 0 => '0') when ps(2)= '1' else     (3 downto 0 => '0') & level2;
   ----------------Synchro barrier, entering cycle 1----------------
   level4<= level3_d1 & (7 downto 0 => '0') when ps_d1(3)= '1' else     (7 downto 0 => '0') & level3_d1;
   R <= level4(28 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                        GenericTable_8_20_F400_uid16
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity GenericTable_8_20_F400_uid16 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          Y : out  std_logic_vector(19 downto 0)   );
end entity;

architecture arch of GenericTable_8_20_F400_uid16 is
signal TableOut :  std_logic_vector(19 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
  with X select TableOut <= 
   "01111111110000010000" when "00000000",
   "01111111010000100000" when "00000001",
   "01111110110000111111" when "00000010",
   "01111110010001101110" when "00000011",
   "01111101110010101100" when "00000100",
   "01111101010011111010" when "00000101",
   "01111100110101010111" when "00000110",
   "01111100010111000010" when "00000111",
   "01111011111000111100" when "00001000",
   "01111011011011000101" when "00001001",
   "01111010111101011100" when "00001010",
   "01111010100000000001" when "00001011",
   "01111010000010110100" when "00001100",
   "01111001100101110101" when "00001101",
   "01111001001001000100" when "00001110",
   "01111000101100100000" when "00001111",
   "01111000010000001010" when "00010000",
   "01110111110100000001" when "00010001",
   "01110111011000000101" when "00010010",
   "01110110111100010110" when "00010011",
   "01110110100000110100" when "00010100",
   "01110110000101011111" when "00010101",
   "01110101101010010110" when "00010110",
   "01110101001111011001" when "00010111",
   "01110100110100101001" when "00011000",
   "01110100011010000110" when "00011001",
   "01110011111111101110" when "00011010",
   "01110011100101100010" when "00011011",
   "01110011001011100001" when "00011100",
   "01110010110001101101" when "00011101",
   "01110010011000000100" when "00011110",
   "01110001111110100110" when "00011111",
   "01110001100101010100" when "00100000",
   "01110001001100001101" when "00100001",
   "01110000110011010001" when "00100010",
   "01110000011010100000" when "00100011",
   "01110000000001111010" when "00100100",
   "01101111101001011110" when "00100101",
   "01101111010001001101" when "00100110",
   "01101110111001000111" when "00100111",
   "01101110100001001011" when "00101000",
   "01101110001001011001" when "00101001",
   "01101101110001110010" when "00101010",
   "01101101011010010100" when "00101011",
   "01101101000011000001" when "00101100",
   "01101100101011110111" when "00101101",
   "01101100010100110111" when "00101110",
   "01101011111110000010" when "00101111",
   "01101011100111010101" when "00110000",
   "01101011010000110010" when "00110001",
   "01101010111010011001" when "00110010",
   "01101010100100001001" when "00110011",
   "01101010001110000010" when "00110100",
   "01101001111000000100" when "00110101",
   "01101001100010001111" when "00110110",
   "01101001001100100011" when "00110111",
   "01101000110111000001" when "00111000",
   "01101000100001100111" when "00111001",
   "01101000001100010101" when "00111010",
   "01100111110111001100" when "00111011",
   "01100111100010001100" when "00111100",
   "01100111001101010101" when "00111101",
   "01100110111000100101" when "00111110",
   "01100110100011111110" when "00111111",
   "01100110001111011111" when "01000000",
   "01100101111011001001" when "01000001",
   "01100101100110111010" when "01000010",
   "01100101010010110011" when "01000011",
   "01100100111110110101" when "01000100",
   "01100100101010111110" when "01000101",
   "01100100010111001111" when "01000110",
   "01100100000011101000" when "01000111",
   "01100011110000001000" when "01001000",
   "01100011011100110000" when "01001001",
   "01100011001001100000" when "01001010",
   "01100010110110010110" when "01001011",
   "01100010100011010101" when "01001100",
   "01100010010000011010" when "01001101",
   "01100001111101100111" when "01001110",
   "01100001101010111011" when "01001111",
   "01100001011000010110" when "01010000",
   "01100001000101111000" when "01010001",
   "01100000110011100001" when "01010010",
   "01100000100001010001" when "01010011",
   "01100000001111001000" when "01010100",
   "01011111111101000110" when "01010101",
   "01011111101011001010" when "01010110",
   "01011111011001010101" when "01010111",
   "01011111000111100111" when "01011000",
   "01011110110110000000" when "01011001",
   "01011110100100011110" when "01011010",
   "01011110010011000011" when "01011011",
   "01011110000001101111" when "01011100",
   "01011101110000100001" when "01011101",
   "01011101011111011001" when "01011110",
   "01011101001110011000" when "01011111",
   "01011100111101011101" when "01100000",
   "01011100101100101000" when "01100001",
   "01011100011011111000" when "01100010",
   "01011100001011001111" when "01100011",
   "01011011111010101100" when "01100100",
   "01011011101010001111" when "01100101",
   "01011011011001111000" when "01100110",
   "01011011001001100110" when "01100111",
   "01011010111001011011" when "01101000",
   "01011010101001010101" when "01101001",
   "01011010011001010100" when "01101010",
   "01011010001001011010" when "01101011",
   "01011001111001100101" when "01101100",
   "01011001101001110101" when "01101101",
   "01011001011010001011" when "01101110",
   "01011001001010100111" when "01101111",
   "01011000111011001000" when "01110000",
   "01011000101011101110" when "01110001",
   "01011000011100011001" when "01110010",
   "01011000001101001010" when "01110011",
   "01010111111110000000" when "01110100",
   "01010111101110111100" when "01110101",
   "01010111011111111100" when "01110110",
   "01010111010001000001" when "01110111",
   "01010111000010001100" when "01111000",
   "01010110110011011100" when "01111001",
   "01010110100100110000" when "01111010",
   "01010110010110001010" when "01111011",
   "01010110000111101000" when "01111100",
   "01010101111001001100" when "01111101",
   "01010101101010110100" when "01111110",
   "01010101011100100001" when "01111111",
   "01010101001110010011" when "10000000",
   "01010101000000001001" when "10000001",
   "01010100110010000100" when "10000010",
   "01010100100100000100" when "10000011",
   "01010100010110001000" when "10000100",
   "01010100001000010001" when "10000101",
   "01010011111010011111" when "10000110",
   "01010011101100110001" when "10000111",
   "01010011011111000111" when "10001000",
   "01010011010001100010" when "10001001",
   "01010011000100000010" when "10001010",
   "01010010110110100101" when "10001011",
   "01010010101001001101" when "10001100",
   "01010010011011111010" when "10001101",
   "01010010001110101010" when "10001110",
   "01010010000001011111" when "10001111",
   "01010001110100011000" when "10010000",
   "01010001100111010110" when "10010001",
   "01010001011010010111" when "10010010",
   "01010001001101011101" when "10010011",
   "01010001000000100110" when "10010100",
   "01010000110011110100" when "10010101",
   "01010000100111000110" when "10010110",
   "01010000011010011011" when "10010111",
   "01010000001101110101" when "10011000",
   "01010000000001010011" when "10011001",
   "01001111110100110100" when "10011010",
   "01001111101000011010" when "10011011",
   "01001111011100000011" when "10011100",
   "01001111001111110000" when "10011101",
   "01001111000011100001" when "10011110",
   "01001110110111010110" when "10011111",
   "01001110101011001110" when "10100000",
   "01001110011111001010" when "10100001",
   "01001110010011001010" when "10100010",
   "01001110000111001101" when "10100011",
   "01001101111011010100" when "10100100",
   "01001101101111011111" when "10100101",
   "01001101100011101101" when "10100110",
   "01001101010111111111" when "10100111",
   "01001101001100010101" when "10101000",
   "01001101000000101110" when "10101001",
   "01001100110101001010" when "10101010",
   "01001100101001101010" when "10101011",
   "01001100011110001101" when "10101100",
   "01001100010010110100" when "10101101",
   "01001100000111011110" when "10101110",
   "01001011111100001011" when "10101111",
   "01001011110000111100" when "10110000",
   "01001011100101110000" when "10110001",
   "01001011011010101000" when "10110010",
   "01001011001111100010" when "10110011",
   "01001011000100100000" when "10110100",
   "01001010111001100001" when "10110101",
   "01001010101110100110" when "10110110",
   "01001010100011101101" when "10110111",
   "01001010011000111000" when "10111000",
   "01001010001110000110" when "10111001",
   "01001010000011010111" when "10111010",
   "01001001111000101011" when "10111011",
   "01001001101110000010" when "10111100",
   "01001001100011011100" when "10111101",
   "01001001011000111001" when "10111110",
   "01001001001110011001" when "10111111",
   "01001001000011111101" when "11000000",
   "01001000111001100011" when "11000001",
   "01001000101111001100" when "11000010",
   "01001000100100111000" when "11000011",
   "01001000011010100111" when "11000100",
   "01001000010000011001" when "11000101",
   "01001000000110001110" when "11000110",
   "01000111111100000110" when "11000111",
   "01000111110010000000" when "11001000",
   "01000111100111111101" when "11001001",
   "01000111011101111110" when "11001010",
   "01000111010100000000" when "11001011",
   "01000111001010000110" when "11001100",
   "01000111000000001111" when "11001101",
   "01000110110110011010" when "11001110",
   "01000110101100101000" when "11001111",
   "01000110100010111000" when "11010000",
   "01000110011001001011" when "11010001",
   "01000110001111100001" when "11010010",
   "01000110000101111010" when "11010011",
   "01000101111100010101" when "11010100",
   "01000101110010110011" when "11010101",
   "01000101101001010011" when "11010110",
   "01000101011111110110" when "11010111",
   "01000101010110011100" when "11011000",
   "01000101001101000100" when "11011001",
   "01000101000011101110" when "11011010",
   "01000100111010011011" when "11011011",
   "01000100110001001011" when "11011100",
   "01000100100111111101" when "11011101",
   "01000100011110110010" when "11011110",
   "01000100010101101001" when "11011111",
   "01000100001100100010" when "11100000",
   "01000100000011011110" when "11100001",
   "01000011111010011100" when "11100010",
   "01000011110001011101" when "11100011",
   "01000011101000100000" when "11100100",
   "01000011011111100101" when "11100101",
   "01000011010110101101" when "11100110",
   "01000011001101110111" when "11100111",
   "01000011000101000100" when "11101000",
   "01000010111100010010" when "11101001",
   "01000010110011100011" when "11101010",
   "01000010101010110110" when "11101011",
   "01000010100010001100" when "11101100",
   "01000010011001100100" when "11101101",
   "01000010010000111110" when "11101110",
   "01000010001000011010" when "11101111",
   "01000001111111111000" when "11110000",
   "01000001110111011001" when "11110001",
   "01000001101110111100" when "11110010",
   "01000001100110100001" when "11110011",
   "01000001011110001000" when "11110100",
   "01000001010101110001" when "11110101",
   "01000001001101011100" when "11110110",
   "01000001000101001010" when "11110111",
   "01000000111100111001" when "11111000",
   "01000000110100101011" when "11111001",
   "01000000101100011111" when "11111010",
   "01000000100100010101" when "11111011",
   "01000000011100001101" when "11111100",
   "01000000010100000111" when "11111101",
   "01000000001100000010" when "11111110",
   "01000000000100000000" when "11111111",
   "--------------------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                        GenericTable_9_12_F400_uid20
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity GenericTable_9_12_F400_uid20 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of GenericTable_9_12_F400_uid20 is
signal TableOut :  std_logic_vector(11 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
  with X select TableOut <= 
   "001110110100" when "000000000",
   "001110010110" when "000000001",
   "001101111000" when "000000010",
   "001101011010" when "000000011",
   "001100111100" when "000000100",
   "001100011101" when "000000101",
   "001011111111" when "000000110",
   "001011100001" when "000000111",
   "001011000011" when "000001000",
   "001010100101" when "000001001",
   "001010000111" when "000001010",
   "001001101001" when "000001011",
   "001001001011" when "000001100",
   "001000101101" when "000001101",
   "001000001111" when "000001110",
   "000111110001" when "000001111",
   "000111010010" when "000010000",
   "000110110100" when "000010001",
   "000110010110" when "000010010",
   "000101111000" when "000010011",
   "000101011010" when "000010100",
   "000100111100" when "000010101",
   "000100011110" when "000010110",
   "000100000000" when "000010111",
   "000011100010" when "000011000",
   "000011000100" when "000011001",
   "000010100110" when "000011010",
   "000010000111" when "000011011",
   "000001101001" when "000011100",
   "000001001011" when "000011101",
   "000000101101" when "000011110",
   "000000001111" when "000011111",
   "001101001011" when "000100000",
   "001100110000" when "000100001",
   "001100010101" when "000100010",
   "001011111010" when "000100011",
   "001011100000" when "000100100",
   "001011000101" when "000100101",
   "001010101010" when "000100110",
   "001010001111" when "000100111",
   "001001110101" when "000101000",
   "001001011010" when "000101001",
   "001000111111" when "000101010",
   "001000100100" when "000101011",
   "001000001010" when "000101100",
   "000111101111" when "000101101",
   "000111010100" when "000101110",
   "000110111001" when "000101111",
   "000110011111" when "000110000",
   "000110000100" when "000110001",
   "000101101001" when "000110010",
   "000101001110" when "000110011",
   "000100110100" when "000110100",
   "000100011001" when "000110101",
   "000011111110" when "000110110",
   "000011100011" when "000110111",
   "000011001001" when "000111000",
   "000010101110" when "000111001",
   "000010010011" when "000111010",
   "000001111000" when "000111011",
   "000001011110" when "000111100",
   "000001000011" when "000111101",
   "000000101000" when "000111110",
   "000000001101" when "000111111",
   "001011110010" when "001000000",
   "001011011010" when "001000001",
   "001011000010" when "001000010",
   "001010101010" when "001000011",
   "001010010010" when "001000100",
   "001001111010" when "001000101",
   "001001100010" when "001000110",
   "001001001010" when "001000111",
   "001000110011" when "001001000",
   "001000011011" when "001001001",
   "001000000011" when "001001010",
   "000111101011" when "001001011",
   "000111010011" when "001001100",
   "000110111011" when "001001101",
   "000110100011" when "001001110",
   "000110001011" when "001001111",
   "000101110011" when "001010000",
   "000101011011" when "001010001",
   "000101000011" when "001010010",
   "000100101011" when "001010011",
   "000100010011" when "001010100",
   "000011111011" when "001010101",
   "000011100011" when "001010110",
   "000011001011" when "001010111",
   "000010110100" when "001011000",
   "000010011100" when "001011001",
   "000010000100" when "001011010",
   "000001101100" when "001011011",
   "000001010100" when "001011100",
   "000000111100" when "001011101",
   "000000100100" when "001011110",
   "000000001100" when "001011111",
   "001010100111" when "001100000",
   "001010010001" when "001100001",
   "001001111100" when "001100010",
   "001001100110" when "001100011",
   "001001010000" when "001100100",
   "001000111011" when "001100101",
   "001000100101" when "001100110",
   "001000010000" when "001100111",
   "000111111010" when "001101000",
   "000111100101" when "001101001",
   "000111001111" when "001101010",
   "000110111010" when "001101011",
   "000110100100" when "001101100",
   "000110001111" when "001101101",
   "000101111001" when "001101110",
   "000101100011" when "001101111",
   "000101001110" when "001110000",
   "000100111000" when "001110001",
   "000100100011" when "001110010",
   "000100001101" when "001110011",
   "000011111000" when "001110100",
   "000011100010" when "001110101",
   "000011001101" when "001110110",
   "000010110111" when "001110111",
   "000010100010" when "001111000",
   "000010001100" when "001111001",
   "000001110110" when "001111010",
   "000001100001" when "001111011",
   "000001001011" when "001111100",
   "000000110110" when "001111101",
   "000000100000" when "001111110",
   "000000001011" when "001111111",
   "001001100110" when "010000000",
   "001001010011" when "010000001",
   "001000111111" when "010000010",
   "001000101100" when "010000011",
   "001000011000" when "010000100",
   "001000000101" when "010000101",
   "000111110001" when "010000110",
   "000111011110" when "010000111",
   "000111001010" when "010001000",
   "000110110111" when "010001001",
   "000110100011" when "010001010",
   "000110010000" when "010001011",
   "000101111100" when "010001100",
   "000101101001" when "010001101",
   "000101010101" when "010001110",
   "000101000010" when "010001111",
   "000100101110" when "010010000",
   "000100011011" when "010010001",
   "000100000111" when "010010010",
   "000011110100" when "010010011",
   "000011100000" when "010010100",
   "000011001101" when "010010101",
   "000010111001" when "010010110",
   "000010100110" when "010010111",
   "000010010010" when "010011000",
   "000001111111" when "010011001",
   "000001101011" when "010011010",
   "000001011000" when "010011011",
   "000001000100" when "010011100",
   "000000110001" when "010011101",
   "000000011101" when "010011110",
   "000000001010" when "010011111",
   "001000101110" when "010100000",
   "001000011101" when "010100001",
   "001000001011" when "010100010",
   "000111111001" when "010100011",
   "000111100111" when "010100100",
   "000111010110" when "010100101",
   "000111000100" when "010100110",
   "000110110010" when "010100111",
   "000110100000" when "010101000",
   "000110001111" when "010101001",
   "000101111101" when "010101010",
   "000101101011" when "010101011",
   "000101011010" when "010101100",
   "000101001000" when "010101101",
   "000100110110" when "010101110",
   "000100100100" when "010101111",
   "000100010011" when "010110000",
   "000100000001" when "010110001",
   "000011101111" when "010110010",
   "000011011110" when "010110011",
   "000011001100" when "010110100",
   "000010111010" when "010110101",
   "000010101000" when "010110110",
   "000010010111" when "010110111",
   "000010000101" when "010111000",
   "000001110011" when "010111001",
   "000001100001" when "010111010",
   "000001010000" when "010111011",
   "000000111110" when "010111100",
   "000000101100" when "010111101",
   "000000011011" when "010111110",
   "000000001001" when "010111111",
   "000111111110" when "011000000",
   "000111101110" when "011000001",
   "000111011101" when "011000010",
   "000111001101" when "011000011",
   "000110111101" when "011000100",
   "000110101101" when "011000101",
   "000110011101" when "011000110",
   "000110001100" when "011000111",
   "000101111100" when "011001000",
   "000101101100" when "011001001",
   "000101011100" when "011001010",
   "000101001100" when "011001011",
   "000100111100" when "011001100",
   "000100101011" when "011001101",
   "000100011011" when "011001110",
   "000100001011" when "011001111",
   "000011111011" when "011010000",
   "000011101011" when "011010001",
   "000011011010" when "011010010",
   "000011001010" when "011010011",
   "000010111010" when "011010100",
   "000010101010" when "011010101",
   "000010011010" when "011010110",
   "000010001010" when "011010111",
   "000001111001" when "011011000",
   "000001101001" when "011011001",
   "000001011001" when "011011010",
   "000001001001" when "011011011",
   "000000111001" when "011011100",
   "000000101000" when "011011101",
   "000000011000" when "011011110",
   "000000001000" when "011011111",
   "000111010011" when "011100000",
   "000111000100" when "011100001",
   "000110110110" when "011100010",
   "000110100111" when "011100011",
   "000110011000" when "011100100",
   "000110001001" when "011100101",
   "000101111010" when "011100110",
   "000101101011" when "011100111",
   "000101011101" when "011101000",
   "000101001110" when "011101001",
   "000100111111" when "011101010",
   "000100110000" when "011101011",
   "000100100001" when "011101100",
   "000100010010" when "011101101",
   "000100000100" when "011101110",
   "000011110101" when "011101111",
   "000011100110" when "011110000",
   "000011010111" when "011110001",
   "000011001000" when "011110010",
   "000010111001" when "011110011",
   "000010101011" when "011110100",
   "000010011100" when "011110101",
   "000010001101" when "011110110",
   "000001111110" when "011110111",
   "000001101111" when "011111000",
   "000001100000" when "011111001",
   "000001010010" when "011111010",
   "000001000011" when "011111011",
   "000000110100" when "011111100",
   "000000100101" when "011111101",
   "000000010110" when "011111110",
   "000000000111" when "011111111",
   "000110101110" when "100000000",
   "000110100000" when "100000001",
   "000110010011" when "100000010",
   "000110000101" when "100000011",
   "000101110111" when "100000100",
   "000101101010" when "100000101",
   "000101011100" when "100000110",
   "000101001110" when "100000111",
   "000101000001" when "100001000",
   "000100110011" when "100001001",
   "000100100101" when "100001010",
   "000100011000" when "100001011",
   "000100001010" when "100001100",
   "000011111100" when "100001101",
   "000011101111" when "100001110",
   "000011100001" when "100001111",
   "000011010100" when "100010000",
   "000011000110" when "100010001",
   "000010111000" when "100010010",
   "000010101011" when "100010011",
   "000010011101" when "100010100",
   "000010001111" when "100010101",
   "000010000010" when "100010110",
   "000001110100" when "100010111",
   "000001100110" when "100011000",
   "000001011001" when "100011001",
   "000001001011" when "100011010",
   "000000111101" when "100011011",
   "000000110000" when "100011100",
   "000000100010" when "100011101",
   "000000010100" when "100011110",
   "000000000111" when "100011111",
   "000110001101" when "100100000",
   "000110000000" when "100100001",
   "000101110100" when "100100010",
   "000101100111" when "100100011",
   "000101011010" when "100100100",
   "000101001110" when "100100101",
   "000101000001" when "100100110",
   "000100110101" when "100100111",
   "000100101000" when "100101000",
   "000100011011" when "100101001",
   "000100001111" when "100101010",
   "000100000010" when "100101011",
   "000011110110" when "100101100",
   "000011101001" when "100101101",
   "000011011100" when "100101110",
   "000011010000" when "100101111",
   "000011000011" when "100110000",
   "000010110111" when "100110001",
   "000010101010" when "100110010",
   "000010011101" when "100110011",
   "000010010001" when "100110100",
   "000010000100" when "100110101",
   "000001111000" when "100110110",
   "000001101011" when "100110111",
   "000001011110" when "100111000",
   "000001010010" when "100111001",
   "000001000101" when "100111010",
   "000000111001" when "100111011",
   "000000101100" when "100111100",
   "000000011111" when "100111101",
   "000000010011" when "100111110",
   "000000000110" when "100111111",
   "000101101111" when "101000000",
   "000101100100" when "101000001",
   "000101011000" when "101000010",
   "000101001100" when "101000011",
   "000101000001" when "101000100",
   "000100110101" when "101000101",
   "000100101001" when "101000110",
   "000100011110" when "101000111",
   "000100010010" when "101001000",
   "000100000110" when "101001001",
   "000011111011" when "101001010",
   "000011101111" when "101001011",
   "000011100011" when "101001100",
   "000011011000" when "101001101",
   "000011001100" when "101001110",
   "000011000000" when "101001111",
   "000010110101" when "101010000",
   "000010101001" when "101010001",
   "000010011101" when "101010010",
   "000010010010" when "101010011",
   "000010000110" when "101010100",
   "000001111010" when "101010101",
   "000001101111" when "101010110",
   "000001100011" when "101010111",
   "000001010111" when "101011000",
   "000001001100" when "101011001",
   "000001000000" when "101011010",
   "000000110100" when "101011011",
   "000000101001" when "101011100",
   "000000011101" when "101011101",
   "000000010001" when "101011110",
   "000000000110" when "101011111",
   "000101010101" when "101100000",
   "000101001010" when "101100001",
   "000101000000" when "101100010",
   "000100110101" when "101100011",
   "000100101010" when "101100100",
   "000100011111" when "101100101",
   "000100010100" when "101100110",
   "000100001001" when "101100111",
   "000011111111" when "101101000",
   "000011110100" when "101101001",
   "000011101001" when "101101010",
   "000011011110" when "101101011",
   "000011010011" when "101101100",
   "000011001000" when "101101101",
   "000010111110" when "101101110",
   "000010110011" when "101101111",
   "000010101000" when "101110000",
   "000010011101" when "101110001",
   "000010010010" when "101110010",
   "000010000111" when "101110011",
   "000001111101" when "101110100",
   "000001110010" when "101110101",
   "000001100111" when "101110110",
   "000001011100" when "101110111",
   "000001010001" when "101111000",
   "000001000110" when "101111001",
   "000000111100" when "101111010",
   "000000110001" when "101111011",
   "000000100110" when "101111100",
   "000000011011" when "101111101",
   "000000010000" when "101111110",
   "000000000101" when "101111111",
   "000100111110" when "110000000",
   "000100110100" when "110000001",
   "000100101010" when "110000010",
   "000100011111" when "110000011",
   "000100010101" when "110000100",
   "000100001011" when "110000101",
   "000100000001" when "110000110",
   "000011110111" when "110000111",
   "000011101101" when "110001000",
   "000011100011" when "110001001",
   "000011011001" when "110001010",
   "000011001111" when "110001011",
   "000011000101" when "110001100",
   "000010111011" when "110001101",
   "000010110001" when "110001110",
   "000010100110" when "110001111",
   "000010011100" when "110010000",
   "000010010010" when "110010001",
   "000010001000" when "110010010",
   "000001111110" when "110010011",
   "000001110100" when "110010100",
   "000001101010" when "110010101",
   "000001100000" when "110010110",
   "000001010110" when "110010111",
   "000001001100" when "110011000",
   "000001000010" when "110011001",
   "000000110111" when "110011010",
   "000000101101" when "110011011",
   "000000100011" when "110011100",
   "000000011001" when "110011101",
   "000000001111" when "110011110",
   "000000000101" when "110011111",
   "000100101001" when "110100000",
   "000100011111" when "110100001",
   "000100010110" when "110100010",
   "000100001100" when "110100011",
   "000100000011" when "110100100",
   "000011111001" when "110100101",
   "000011110000" when "110100110",
   "000011100111" when "110100111",
   "000011011101" when "110101000",
   "000011010100" when "110101001",
   "000011001010" when "110101010",
   "000011000001" when "110101011",
   "000010111000" when "110101100",
   "000010101110" when "110101101",
   "000010100101" when "110101110",
   "000010011011" when "110101111",
   "000010010010" when "110110000",
   "000010001000" when "110110001",
   "000001111111" when "110110010",
   "000001110110" when "110110011",
   "000001101100" when "110110100",
   "000001100011" when "110110101",
   "000001011001" when "110110110",
   "000001010000" when "110110111",
   "000001000111" when "110111000",
   "000000111101" when "110111001",
   "000000110100" when "110111010",
   "000000101010" when "110111011",
   "000000100001" when "110111100",
   "000000011000" when "110111101",
   "000000001110" when "110111110",
   "000000000101" when "110111111",
   "000100010101" when "111000000",
   "000100001101" when "111000001",
   "000100000100" when "111000010",
   "000011111011" when "111000011",
   "000011110010" when "111000100",
   "000011101001" when "111000101",
   "000011100001" when "111000110",
   "000011011000" when "111000111",
   "000011001111" when "111001000",
   "000011000110" when "111001001",
   "000010111101" when "111001010",
   "000010110101" when "111001011",
   "000010101100" when "111001100",
   "000010100011" when "111001101",
   "000010011010" when "111001110",
   "000010010001" when "111001111",
   "000010001001" when "111010000",
   "000010000000" when "111010001",
   "000001110111" when "111010010",
   "000001101110" when "111010011",
   "000001100101" when "111010100",
   "000001011100" when "111010101",
   "000001010100" when "111010110",
   "000001001011" when "111010111",
   "000001000010" when "111011000",
   "000000111001" when "111011001",
   "000000110000" when "111011010",
   "000000101000" when "111011011",
   "000000011111" when "111011100",
   "000000010110" when "111011101",
   "000000001101" when "111011110",
   "000000000100" when "111011111",
   "000100000100" when "111100000",
   "000011111100" when "111100001",
   "000011110100" when "111100010",
   "000011101011" when "111100011",
   "000011100011" when "111100100",
   "000011011011" when "111100101",
   "000011010011" when "111100110",
   "000011001010" when "111100111",
   "000011000010" when "111101000",
   "000010111010" when "111101001",
   "000010110010" when "111101010",
   "000010101001" when "111101011",
   "000010100001" when "111101100",
   "000010011001" when "111101101",
   "000010010000" when "111101110",
   "000010001000" when "111101111",
   "000010000000" when "111110000",
   "000001111000" when "111110001",
   "000001101111" when "111110010",
   "000001100111" when "111110011",
   "000001011111" when "111110100",
   "000001010111" when "111110101",
   "000001001110" when "111110110",
   "000001000110" when "111110111",
   "000000111110" when "111111000",
   "000000110110" when "111111001",
   "000000101101" when "111111010",
   "000000100101" when "111111011",
   "000000011101" when "111111100",
   "000000010101" when "111111101",
   "000000001100" when "111111110",
   "000000000100" when "111111111",
   "------------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                              reciprocal_uid23
--        (BipartiteTable_f_2_1Px_M1bM16_in_M14_out_1_M16_F400_uid14)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Matei Istoan (2014)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity reciprocal_uid23 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(13 downto 0);
          Y : out  std_logic_vector(17 downto 0)   );
end entity;

architecture arch of reciprocal_uid23 is
   component GenericTable_8_20_F400_uid16 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             Y : out  std_logic_vector(19 downto 0)   );
   end component;

   component GenericTable_9_12_F400_uid20 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(11 downto 0)   );
   end component;

signal X0 :  std_logic_vector(3 downto 0);
signal X1 :  std_logic_vector(3 downto 0);
signal X2 :  std_logic_vector(5 downto 0);
signal X2_msb :  std_logic;
signal X2_short :  std_logic_vector(4 downto 0);
signal X2_short_inv :  std_logic_vector(4 downto 0);
signal tableTIVaddr :  std_logic_vector(7 downto 0);
signal tableTOaddr :  std_logic_vector(8 downto 0);
signal tableTIVout :  std_logic_vector(19 downto 0);
signal tableTOout :  std_logic_vector(11 downto 0);
signal tableTOout_inv :  std_logic_vector(11 downto 0);
signal tableTIV_fxp :  signed(1+18 downto 0);
signal tableTO_fxp :  signed(-7+18 downto 0);
signal tableTO_fxp_sgnExt :  signed(1+18 downto 0);
signal Y_int :  signed(1+18 downto 0);
signal Y_int_short :  signed(1+17 downto 0);
signal Y_rnd :  signed(1+17 downto 0);
attribute rom_extract: string;
attribute rom_style: string;
attribute rom_extract of GenericTable_8_20_F400_uid16: component is "yes";
attribute rom_extract of GenericTable_9_12_F400_uid20: component is "yes";
attribute rom_style of GenericTable_8_20_F400_uid16: component is "block";
attribute rom_style of GenericTable_9_12_F400_uid20: component is "block";
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   X0 <= X(13 downto 10);
   X1 <= X(9 downto 6);
   X2 <= X(5 downto 0);

   X2_msb <= X2(5);
   X2_short <= X2(4 downto 0);
   X2_short_inv <= X2_short xor (4 downto 0 => X2_msb);

   tableTIVaddr <= X0 & X1;
   tableTOaddr <= X0 & X2_short_inv;

   TIVtable: GenericTable_8_20_F400_uid16  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => tableTIVaddr,
                 Y => tableTIVout);

   TOtable: GenericTable_9_12_F400_uid20  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => tableTOaddr,
                 Y => tableTOout);

   tableTOout_inv <= tableTOout xor (11 downto 0 => X2_msb);

   tableTIV_fxp <= signed(tableTIVout);
   tableTO_fxp <= signed(tableTOout_inv);
   tableTO_fxp_sgnExt <= (7 downto 0 => tableTO_fxp(11)) & tableTO_fxp(11 downto 0); -- fix resize from (-7, -18) to (1, -18)

   Y_int <= tableTIV_fxp + tableTO_fxp_sgnExt;
   Y_int_short <= Y_int(19 downto 1); -- fix resize from (1, -18) to (1, -17)
   Y_rnd <= Y_int_short + ("000000000000000000" & '1');
   Y <= std_logic_vector(Y_rnd(18 downto 1));
end architecture;

--------------------------------------------------------------------------------
--                       GenericTable_10_16_F400_uid29
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity GenericTable_10_16_F400_uid29 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(15 downto 0)   );
end entity;

architecture arch of GenericTable_10_16_F400_uid29 is
signal TableOut, TableOut_d1 :  std_logic_vector(15 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            TableOut_d1 <=  TableOut;
         end if;
      end process;
  with X select TableOut <= 
   "0000000000010100" when "0000000000",
   "0000000000111101" when "0000000001",
   "0000000001100110" when "0000000010",
   "0000000010001110" when "0000000011",
   "0000000010110111" when "0000000100",
   "0000000011100000" when "0000000101",
   "0000000100001001" when "0000000110",
   "0000000100110001" when "0000000111",
   "0000000101011010" when "0000001000",
   "0000000110000011" when "0000001001",
   "0000000110101011" when "0000001010",
   "0000000111010100" when "0000001011",
   "0000000111111101" when "0000001100",
   "0000001000100110" when "0000001101",
   "0000001001001110" when "0000001110",
   "0000001001110111" when "0000001111",
   "0000001010100000" when "0000010000",
   "0000001011001001" when "0000010001",
   "0000001011110001" when "0000010010",
   "0000001100011010" when "0000010011",
   "0000001101000011" when "0000010100",
   "0000001101101100" when "0000010101",
   "0000001110010100" when "0000010110",
   "0000001110111101" when "0000010111",
   "0000001111100110" when "0000011000",
   "0000010000001110" when "0000011001",
   "0000010000110111" when "0000011010",
   "0000010001100000" when "0000011011",
   "0000010010001001" when "0000011100",
   "0000010010110001" when "0000011101",
   "0000010011011010" when "0000011110",
   "0000010100000011" when "0000011111",
   "0000010100101011" when "0000100000",
   "0000010101010100" when "0000100001",
   "0000010101111101" when "0000100010",
   "0000010110100110" when "0000100011",
   "0000010111001110" when "0000100100",
   "0000010111110111" when "0000100101",
   "0000011000100000" when "0000100110",
   "0000011001001000" when "0000100111",
   "0000011001110001" when "0000101000",
   "0000011010011010" when "0000101001",
   "0000011011000010" when "0000101010",
   "0000011011101011" when "0000101011",
   "0000011100010100" when "0000101100",
   "0000011100111100" when "0000101101",
   "0000011101100101" when "0000101110",
   "0000011110001110" when "0000101111",
   "0000011110110110" when "0000110000",
   "0000011111011111" when "0000110001",
   "0000100000001000" when "0000110010",
   "0000100000110000" when "0000110011",
   "0000100001011001" when "0000110100",
   "0000100010000001" when "0000110101",
   "0000100010101010" when "0000110110",
   "0000100011010011" when "0000110111",
   "0000100011111011" when "0000111000",
   "0000100100100100" when "0000111001",
   "0000100101001101" when "0000111010",
   "0000100101110101" when "0000111011",
   "0000100110011110" when "0000111100",
   "0000100111000110" when "0000111101",
   "0000100111101111" when "0000111110",
   "0000101000011000" when "0000111111",
   "0000101001000000" when "0001000000",
   "0000101001101001" when "0001000001",
   "0000101010010001" when "0001000010",
   "0000101010111010" when "0001000011",
   "0000101011100010" when "0001000100",
   "0000101100001011" when "0001000101",
   "0000101100110100" when "0001000110",
   "0000101101011100" when "0001000111",
   "0000101110000101" when "0001001000",
   "0000101110101101" when "0001001001",
   "0000101111010110" when "0001001010",
   "0000101111111110" when "0001001011",
   "0000110000100111" when "0001001100",
   "0000110001001111" when "0001001101",
   "0000110001111000" when "0001001110",
   "0000110010100000" when "0001001111",
   "0000110011001001" when "0001010000",
   "0000110011110001" when "0001010001",
   "0000110100011010" when "0001010010",
   "0000110101000010" when "0001010011",
   "0000110101101011" when "0001010100",
   "0000110110010011" when "0001010101",
   "0000110110111100" when "0001010110",
   "0000110111100100" when "0001010111",
   "0000111000001101" when "0001011000",
   "0000111000110101" when "0001011001",
   "0000111001011101" when "0001011010",
   "0000111010000110" when "0001011011",
   "0000111010101110" when "0001011100",
   "0000111011010111" when "0001011101",
   "0000111011111111" when "0001011110",
   "0000111100100111" when "0001011111",
   "0000111101010000" when "0001100000",
   "0000111101111000" when "0001100001",
   "0000111110100001" when "0001100010",
   "0000111111001001" when "0001100011",
   "0000111111110001" when "0001100100",
   "0001000000011010" when "0001100101",
   "0001000001000010" when "0001100110",
   "0001000001101010" when "0001100111",
   "0001000010010011" when "0001101000",
   "0001000010111011" when "0001101001",
   "0001000011100011" when "0001101010",
   "0001000100001100" when "0001101011",
   "0001000100110100" when "0001101100",
   "0001000101011100" when "0001101101",
   "0001000110000101" when "0001101110",
   "0001000110101101" when "0001101111",
   "0001000111010101" when "0001110000",
   "0001000111111101" when "0001110001",
   "0001001000100110" when "0001110010",
   "0001001001001110" when "0001110011",
   "0001001001110110" when "0001110100",
   "0001001010011110" when "0001110101",
   "0001001011000110" when "0001110110",
   "0001001011101111" when "0001110111",
   "0001001100010111" when "0001111000",
   "0001001100111111" when "0001111001",
   "0001001101100111" when "0001111010",
   "0001001110001111" when "0001111011",
   "0001001110111000" when "0001111100",
   "0001001111100000" when "0001111101",
   "0001010000001000" when "0001111110",
   "0001010000110000" when "0001111111",
   "0001010001011000" when "0010000000",
   "0001010010000000" when "0010000001",
   "0001010010101000" when "0010000010",
   "0001010011010000" when "0010000011",
   "0001010011111000" when "0010000100",
   "0001010100100000" when "0010000101",
   "0001010101001001" when "0010000110",
   "0001010101110001" when "0010000111",
   "0001010110011001" when "0010001000",
   "0001010111000001" when "0010001001",
   "0001010111101001" when "0010001010",
   "0001011000010001" when "0010001011",
   "0001011000111001" when "0010001100",
   "0001011001100001" when "0010001101",
   "0001011010001001" when "0010001110",
   "0001011010110001" when "0010001111",
   "0001011011011001" when "0010010000",
   "0001011100000000" when "0010010001",
   "0001011100101000" when "0010010010",
   "0001011101010000" when "0010010011",
   "0001011101111000" when "0010010100",
   "0001011110100000" when "0010010101",
   "0001011111001000" when "0010010110",
   "0001011111110000" when "0010010111",
   "0001100000011000" when "0010011000",
   "0001100001000000" when "0010011001",
   "0001100001100111" when "0010011010",
   "0001100010001111" when "0010011011",
   "0001100010110111" when "0010011100",
   "0001100011011111" when "0010011101",
   "0001100100000111" when "0010011110",
   "0001100100101110" when "0010011111",
   "0001100101010110" when "0010100000",
   "0001100101111110" when "0010100001",
   "0001100110100110" when "0010100010",
   "0001100111001110" when "0010100011",
   "0001100111110101" when "0010100100",
   "0001101000011101" when "0010100101",
   "0001101001000101" when "0010100110",
   "0001101001101100" when "0010100111",
   "0001101010010100" when "0010101000",
   "0001101010111100" when "0010101001",
   "0001101011100011" when "0010101010",
   "0001101100001011" when "0010101011",
   "0001101100110011" when "0010101100",
   "0001101101011010" when "0010101101",
   "0001101110000010" when "0010101110",
   "0001101110101001" when "0010101111",
   "0001101111010001" when "0010110000",
   "0001101111111001" when "0010110001",
   "0001110000100000" when "0010110010",
   "0001110001001000" when "0010110011",
   "0001110001101111" when "0010110100",
   "0001110010010111" when "0010110101",
   "0001110010111110" when "0010110110",
   "0001110011100110" when "0010110111",
   "0001110100001101" when "0010111000",
   "0001110100110101" when "0010111001",
   "0001110101011100" when "0010111010",
   "0001110110000011" when "0010111011",
   "0001110110101011" when "0010111100",
   "0001110111010010" when "0010111101",
   "0001110111111010" when "0010111110",
   "0001111000100001" when "0010111111",
   "0001111001001000" when "0011000000",
   "0001111001110000" when "0011000001",
   "0001111010010111" when "0011000010",
   "0001111010111110" when "0011000011",
   "0001111011100110" when "0011000100",
   "0001111100001101" when "0011000101",
   "0001111100110100" when "0011000110",
   "0001111101011011" when "0011000111",
   "0001111110000011" when "0011001000",
   "0001111110101010" when "0011001001",
   "0001111111010001" when "0011001010",
   "0001111111111000" when "0011001011",
   "0010000000100000" when "0011001100",
   "0010000001000111" when "0011001101",
   "0010000001101110" when "0011001110",
   "0010000010010101" when "0011001111",
   "0010000010111100" when "0011010000",
   "0010000011100011" when "0011010001",
   "0010000100001010" when "0011010010",
   "0010000100110001" when "0011010011",
   "0010000101011001" when "0011010100",
   "0010000110000000" when "0011010101",
   "0010000110100111" when "0011010110",
   "0010000111001110" when "0011010111",
   "0010000111110101" when "0011011000",
   "0010001000011100" when "0011011001",
   "0010001001000011" when "0011011010",
   "0010001001101010" when "0011011011",
   "0010001010010001" when "0011011100",
   "0010001010110111" when "0011011101",
   "0010001011011110" when "0011011110",
   "0010001100000101" when "0011011111",
   "0010001100101100" when "0011100000",
   "0010001101010011" when "0011100001",
   "0010001101111010" when "0011100010",
   "0010001110100001" when "0011100011",
   "0010001111001000" when "0011100100",
   "0010001111101110" when "0011100101",
   "0010010000010101" when "0011100110",
   "0010010000111100" when "0011100111",
   "0010010001100011" when "0011101000",
   "0010010010001001" when "0011101001",
   "0010010010110000" when "0011101010",
   "0010010011010111" when "0011101011",
   "0010010011111110" when "0011101100",
   "0010010100100100" when "0011101101",
   "0010010101001011" when "0011101110",
   "0010010101110001" when "0011101111",
   "0010010110011000" when "0011110000",
   "0010010110111111" when "0011110001",
   "0010010111100101" when "0011110010",
   "0010011000001100" when "0011110011",
   "0010011000110010" when "0011110100",
   "0010011001011001" when "0011110101",
   "0010011001111111" when "0011110110",
   "0010011010100110" when "0011110111",
   "0010011011001100" when "0011111000",
   "0010011011110011" when "0011111001",
   "0010011100011001" when "0011111010",
   "0010011101000000" when "0011111011",
   "0010011101100110" when "0011111100",
   "0010011110001101" when "0011111101",
   "0010011110110011" when "0011111110",
   "0010011111011001" when "0011111111",
   "0010100000000000" when "0100000000",
   "0010100000100110" when "0100000001",
   "0010100001001100" when "0100000010",
   "0010100001110011" when "0100000011",
   "0010100010011001" when "0100000100",
   "0010100010111111" when "0100000101",
   "0010100011100101" when "0100000110",
   "0010100100001100" when "0100000111",
   "0010100100110010" when "0100001000",
   "0010100101011000" when "0100001001",
   "0010100101111110" when "0100001010",
   "0010100110100100" when "0100001011",
   "0010100111001011" when "0100001100",
   "0010100111110001" when "0100001101",
   "0010101000010111" when "0100001110",
   "0010101000111101" when "0100001111",
   "0010101001100011" when "0100010000",
   "0010101010001001" when "0100010001",
   "0010101010101111" when "0100010010",
   "0010101011010101" when "0100010011",
   "0010101011111011" when "0100010100",
   "0010101100100001" when "0100010101",
   "0010101101000111" when "0100010110",
   "0010101101101101" when "0100010111",
   "0010101110010011" when "0100011000",
   "0010101110111001" when "0100011001",
   "0010101111011110" when "0100011010",
   "0010110000000100" when "0100011011",
   "0010110000101010" when "0100011100",
   "0010110001010000" when "0100011101",
   "0010110001110110" when "0100011110",
   "0010110010011011" when "0100011111",
   "0010110011000001" when "0100100000",
   "0010110011100111" when "0100100001",
   "0010110100001101" when "0100100010",
   "0010110100110010" when "0100100011",
   "0010110101011000" when "0100100100",
   "0010110101111110" when "0100100101",
   "0010110110100011" when "0100100110",
   "0010110111001001" when "0100100111",
   "0010110111101111" when "0100101000",
   "0010111000010100" when "0100101001",
   "0010111000111010" when "0100101010",
   "0010111001011111" when "0100101011",
   "0010111010000101" when "0100101100",
   "0010111010101010" when "0100101101",
   "0010111011010000" when "0100101110",
   "0010111011110101" when "0100101111",
   "0010111100011011" when "0100110000",
   "0010111101000000" when "0100110001",
   "0010111101100110" when "0100110010",
   "0010111110001011" when "0100110011",
   "0010111110110000" when "0100110100",
   "0010111111010110" when "0100110101",
   "0010111111111011" when "0100110110",
   "0011000000100000" when "0100110111",
   "0011000001000110" when "0100111000",
   "0011000001101011" when "0100111001",
   "0011000010010000" when "0100111010",
   "0011000010110101" when "0100111011",
   "0011000011011010" when "0100111100",
   "0011000100000000" when "0100111101",
   "0011000100100101" when "0100111110",
   "0011000101001010" when "0100111111",
   "0011000101101111" when "0101000000",
   "0011000110010100" when "0101000001",
   "0011000110111001" when "0101000010",
   "0011000111011110" when "0101000011",
   "0011001000000011" when "0101000100",
   "0011001000101000" when "0101000101",
   "0011001001001101" when "0101000110",
   "0011001001110010" when "0101000111",
   "0011001010010111" when "0101001000",
   "0011001010111100" when "0101001001",
   "0011001011100001" when "0101001010",
   "0011001100000110" when "0101001011",
   "0011001100101011" when "0101001100",
   "0011001101010000" when "0101001101",
   "0011001101110101" when "0101001110",
   "0011001110011001" when "0101001111",
   "0011001110111110" when "0101010000",
   "0011001111100011" when "0101010001",
   "0011010000001000" when "0101010010",
   "0011010000101100" when "0101010011",
   "0011010001010001" when "0101010100",
   "0011010001110110" when "0101010101",
   "0011010010011010" when "0101010110",
   "0011010010111111" when "0101010111",
   "0011010011100100" when "0101011000",
   "0011010100001000" when "0101011001",
   "0011010100101101" when "0101011010",
   "0011010101010001" when "0101011011",
   "0011010101110110" when "0101011100",
   "0011010110011010" when "0101011101",
   "0011010110111111" when "0101011110",
   "0011010111100011" when "0101011111",
   "0011011000001000" when "0101100000",
   "0011011000101100" when "0101100001",
   "0011011001010001" when "0101100010",
   "0011011001110101" when "0101100011",
   "0011011010011001" when "0101100100",
   "0011011010111110" when "0101100101",
   "0011011011100010" when "0101100110",
   "0011011100000110" when "0101100111",
   "0011011100101010" when "0101101000",
   "0011011101001111" when "0101101001",
   "0011011101110011" when "0101101010",
   "0011011110010111" when "0101101011",
   "0011011110111011" when "0101101100",
   "0011011111011111" when "0101101101",
   "0011100000000100" when "0101101110",
   "0011100000101000" when "0101101111",
   "0011100001001100" when "0101110000",
   "0011100001110000" when "0101110001",
   "0011100010010100" when "0101110010",
   "0011100010111000" when "0101110011",
   "0011100011011100" when "0101110100",
   "0011100100000000" when "0101110101",
   "0011100100100100" when "0101110110",
   "0011100101001000" when "0101110111",
   "0011100101101100" when "0101111000",
   "0011100110001111" when "0101111001",
   "0011100110110011" when "0101111010",
   "0011100111010111" when "0101111011",
   "0011100111111011" when "0101111100",
   "0011101000011111" when "0101111101",
   "0011101001000011" when "0101111110",
   "0011101001100110" when "0101111111",
   "0011101010001010" when "0110000000",
   "0011101010101110" when "0110000001",
   "0011101011010001" when "0110000010",
   "0011101011110101" when "0110000011",
   "0011101100011001" when "0110000100",
   "0011101100111100" when "0110000101",
   "0011101101100000" when "0110000110",
   "0011101110000011" when "0110000111",
   "0011101110100111" when "0110001000",
   "0011101111001010" when "0110001001",
   "0011101111101110" when "0110001010",
   "0011110000010001" when "0110001011",
   "0011110000110101" when "0110001100",
   "0011110001011000" when "0110001101",
   "0011110001111100" when "0110001110",
   "0011110010011111" when "0110001111",
   "0011110011000010" when "0110010000",
   "0011110011100110" when "0110010001",
   "0011110100001001" when "0110010010",
   "0011110100101100" when "0110010011",
   "0011110101010000" when "0110010100",
   "0011110101110011" when "0110010101",
   "0011110110010110" when "0110010110",
   "0011110110111001" when "0110010111",
   "0011110111011100" when "0110011000",
   "0011111000000000" when "0110011001",
   "0011111000100011" when "0110011010",
   "0011111001000110" when "0110011011",
   "0011111001101001" when "0110011100",
   "0011111010001100" when "0110011101",
   "0011111010101111" when "0110011110",
   "0011111011010010" when "0110011111",
   "0011111011110101" when "0110100000",
   "0011111100011000" when "0110100001",
   "0011111100111011" when "0110100010",
   "0011111101011110" when "0110100011",
   "0011111110000000" when "0110100100",
   "0011111110100011" when "0110100101",
   "0011111111000110" when "0110100110",
   "0011111111101001" when "0110100111",
   "0100000000001100" when "0110101000",
   "0100000000101110" when "0110101001",
   "0100000001010001" when "0110101010",
   "0100000001110100" when "0110101011",
   "0100000010010111" when "0110101100",
   "0100000010111001" when "0110101101",
   "0100000011011100" when "0110101110",
   "0100000011111111" when "0110101111",
   "0100000100100001" when "0110110000",
   "0100000101000100" when "0110110001",
   "0100000101100110" when "0110110010",
   "0100000110001001" when "0110110011",
   "0100000110101011" when "0110110100",
   "0100000111001110" when "0110110101",
   "0100000111110000" when "0110110110",
   "0100001000010011" when "0110110111",
   "0100001000110101" when "0110111000",
   "0100001001010111" when "0110111001",
   "0100001001111010" when "0110111010",
   "0100001010011100" when "0110111011",
   "0100001010111110" when "0110111100",
   "0100001011100001" when "0110111101",
   "0100001100000011" when "0110111110",
   "0100001100100101" when "0110111111",
   "0100001101000111" when "0111000000",
   "0100001101101001" when "0111000001",
   "0100001110001100" when "0111000010",
   "0100001110101110" when "0111000011",
   "0100001111010000" when "0111000100",
   "0100001111110010" when "0111000101",
   "0100010000010100" when "0111000110",
   "0100010000110110" when "0111000111",
   "0100010001011000" when "0111001000",
   "0100010001111010" when "0111001001",
   "0100010010011100" when "0111001010",
   "0100010010111110" when "0111001011",
   "0100010011100000" when "0111001100",
   "0100010100000010" when "0111001101",
   "0100010100100011" when "0111001110",
   "0100010101000101" when "0111001111",
   "0100010101100111" when "0111010000",
   "0100010110001001" when "0111010001",
   "0100010110101011" when "0111010010",
   "0100010111001100" when "0111010011",
   "0100010111101110" when "0111010100",
   "0100011000010000" when "0111010101",
   "0100011000110001" when "0111010110",
   "0100011001010011" when "0111010111",
   "0100011001110101" when "0111011000",
   "0100011010010110" when "0111011001",
   "0100011010111000" when "0111011010",
   "0100011011011001" when "0111011011",
   "0100011011111011" when "0111011100",
   "0100011100011100" when "0111011101",
   "0100011100111110" when "0111011110",
   "0100011101011111" when "0111011111",
   "0100011110000000" when "0111100000",
   "0100011110100010" when "0111100001",
   "0100011111000011" when "0111100010",
   "0100011111100101" when "0111100011",
   "0100100000000110" when "0111100100",
   "0100100000100111" when "0111100101",
   "0100100001001000" when "0111100110",
   "0100100001101010" when "0111100111",
   "0100100010001011" when "0111101000",
   "0100100010101100" when "0111101001",
   "0100100011001101" when "0111101010",
   "0100100011101110" when "0111101011",
   "0100100100001111" when "0111101100",
   "0100100100110000" when "0111101101",
   "0100100101010010" when "0111101110",
   "0100100101110011" when "0111101111",
   "0100100110010100" when "0111110000",
   "0100100110110101" when "0111110001",
   "0100100111010101" when "0111110010",
   "0100100111110110" when "0111110011",
   "0100101000010111" when "0111110100",
   "0100101000111000" when "0111110101",
   "0100101001011001" when "0111110110",
   "0100101001111010" when "0111110111",
   "0100101010011011" when "0111111000",
   "0100101010111011" when "0111111001",
   "0100101011011100" when "0111111010",
   "0100101011111101" when "0111111011",
   "0100101100011110" when "0111111100",
   "0100101100111110" when "0111111101",
   "0100101101011111" when "0111111110",
   "0100101110000000" when "0111111111",
   "0100101110100000" when "1000000000",
   "0100101111000001" when "1000000001",
   "0100101111100001" when "1000000010",
   "0100110000000010" when "1000000011",
   "0100110000100010" when "1000000100",
   "0100110001000011" when "1000000101",
   "0100110001100011" when "1000000110",
   "0100110010000100" when "1000000111",
   "0100110010100100" when "1000001000",
   "0100110011000100" when "1000001001",
   "0100110011100101" when "1000001010",
   "0100110100000101" when "1000001011",
   "0100110100100101" when "1000001100",
   "0100110101000110" when "1000001101",
   "0100110101100110" when "1000001110",
   "0100110110000110" when "1000001111",
   "0100110110100110" when "1000010000",
   "0100110111000110" when "1000010001",
   "0100110111100110" when "1000010010",
   "0100111000000111" when "1000010011",
   "0100111000100111" when "1000010100",
   "0100111001000111" when "1000010101",
   "0100111001100111" when "1000010110",
   "0100111010000111" when "1000010111",
   "0100111010100111" when "1000011000",
   "0100111011000111" when "1000011001",
   "0100111011100111" when "1000011010",
   "0100111100000111" when "1000011011",
   "0100111100100110" when "1000011100",
   "0100111101000110" when "1000011101",
   "0100111101100110" when "1000011110",
   "0100111110000110" when "1000011111",
   "0100111110100110" when "1000100000",
   "0100111111000101" when "1000100001",
   "0100111111100101" when "1000100010",
   "0101000000000101" when "1000100011",
   "0101000000100101" when "1000100100",
   "0101000001000100" when "1000100101",
   "0101000001100100" when "1000100110",
   "0101000010000011" when "1000100111",
   "0101000010100011" when "1000101000",
   "0101000011000010" when "1000101001",
   "0101000011100010" when "1000101010",
   "0101000100000001" when "1000101011",
   "0101000100100001" when "1000101100",
   "0101000101000000" when "1000101101",
   "0101000101100000" when "1000101110",
   "0101000101111111" when "1000101111",
   "0101000110011111" when "1000110000",
   "0101000110111110" when "1000110001",
   "0101000111011101" when "1000110010",
   "0101000111111101" when "1000110011",
   "0101001000011100" when "1000110100",
   "0101001000111011" when "1000110101",
   "0101001001011010" when "1000110110",
   "0101001001111001" when "1000110111",
   "0101001010011001" when "1000111000",
   "0101001010111000" when "1000111001",
   "0101001011010111" when "1000111010",
   "0101001011110110" when "1000111011",
   "0101001100010101" when "1000111100",
   "0101001100110100" when "1000111101",
   "0101001101010011" when "1000111110",
   "0101001101110010" when "1000111111",
   "0101001110010001" when "1001000000",
   "0101001110110000" when "1001000001",
   "0101001111001111" when "1001000010",
   "0101001111101110" when "1001000011",
   "0101010000001100" when "1001000100",
   "0101010000101011" when "1001000101",
   "0101010001001010" when "1001000110",
   "0101010001101001" when "1001000111",
   "0101010010001000" when "1001001000",
   "0101010010100110" when "1001001001",
   "0101010011000101" when "1001001010",
   "0101010011100100" when "1001001011",
   "0101010100000010" when "1001001100",
   "0101010100100001" when "1001001101",
   "0101010100111111" when "1001001110",
   "0101010101011110" when "1001001111",
   "0101010101111101" when "1001010000",
   "0101010110011011" when "1001010001",
   "0101010110111010" when "1001010010",
   "0101010111011000" when "1001010011",
   "0101010111110110" when "1001010100",
   "0101011000010101" when "1001010101",
   "0101011000110011" when "1001010110",
   "0101011001010010" when "1001010111",
   "0101011001110000" when "1001011000",
   "0101011010001110" when "1001011001",
   "0101011010101101" when "1001011010",
   "0101011011001011" when "1001011011",
   "0101011011101001" when "1001011100",
   "0101011100000111" when "1001011101",
   "0101011100100101" when "1001011110",
   "0101011101000100" when "1001011111",
   "0101011101100010" when "1001100000",
   "0101011110000000" when "1001100001",
   "0101011110011110" when "1001100010",
   "0101011110111100" when "1001100011",
   "0101011111011010" when "1001100100",
   "0101011111111000" when "1001100101",
   "0101100000010110" when "1001100110",
   "0101100000110100" when "1001100111",
   "0101100001010010" when "1001101000",
   "0101100001110000" when "1001101001",
   "0101100010001110" when "1001101010",
   "0101100010101011" when "1001101011",
   "0101100011001001" when "1001101100",
   "0101100011100111" when "1001101101",
   "0101100100000101" when "1001101110",
   "0101100100100010" when "1001101111",
   "0101100101000000" when "1001110000",
   "0101100101011110" when "1001110001",
   "0101100101111011" when "1001110010",
   "0101100110011001" when "1001110011",
   "0101100110110111" when "1001110100",
   "0101100111010100" when "1001110101",
   "0101100111110010" when "1001110110",
   "0101101000001111" when "1001110111",
   "0101101000101101" when "1001111000",
   "0101101001001010" when "1001111001",
   "0101101001101000" when "1001111010",
   "0101101010000101" when "1001111011",
   "0101101010100011" when "1001111100",
   "0101101011000000" when "1001111101",
   "0101101011011101" when "1001111110",
   "0101101011111011" when "1001111111",
   "0101101100011000" when "1010000000",
   "0101101100110101" when "1010000001",
   "0101101101010011" when "1010000010",
   "0101101101110000" when "1010000011",
   "0101101110001101" when "1010000100",
   "0101101110101010" when "1010000101",
   "0101101111000111" when "1010000110",
   "0101101111100100" when "1010000111",
   "0101110000000001" when "1010001000",
   "0101110000011111" when "1010001001",
   "0101110000111100" when "1010001010",
   "0101110001011001" when "1010001011",
   "0101110001110110" when "1010001100",
   "0101110010010011" when "1010001101",
   "0101110010110000" when "1010001110",
   "0101110011001100" when "1010001111",
   "0101110011101001" when "1010010000",
   "0101110100000110" when "1010010001",
   "0101110100100011" when "1010010010",
   "0101110101000000" when "1010010011",
   "0101110101011101" when "1010010100",
   "0101110101111001" when "1010010101",
   "0101110110010110" when "1010010110",
   "0101110110110011" when "1010010111",
   "0101110111010000" when "1010011000",
   "0101110111101100" when "1010011001",
   "0101111000001001" when "1010011010",
   "0101111000100101" when "1010011011",
   "0101111001000010" when "1010011100",
   "0101111001011111" when "1010011101",
   "0101111001111011" when "1010011110",
   "0101111010011000" when "1010011111",
   "0101111010110100" when "1010100000",
   "0101111011010001" when "1010100001",
   "0101111011101101" when "1010100010",
   "0101111100001001" when "1010100011",
   "0101111100100110" when "1010100100",
   "0101111101000010" when "1010100101",
   "0101111101011110" when "1010100110",
   "0101111101111011" when "1010100111",
   "0101111110010111" when "1010101000",
   "0101111110110011" when "1010101001",
   "0101111111001111" when "1010101010",
   "0101111111101100" when "1010101011",
   "0110000000001000" when "1010101100",
   "0110000000100100" when "1010101101",
   "0110000001000000" when "1010101110",
   "0110000001011100" when "1010101111",
   "0110000001111000" when "1010110000",
   "0110000010010100" when "1010110001",
   "0110000010110000" when "1010110010",
   "0110000011001100" when "1010110011",
   "0110000011101000" when "1010110100",
   "0110000100000100" when "1010110101",
   "0110000100100000" when "1010110110",
   "0110000100111100" when "1010110111",
   "0110000101011000" when "1010111000",
   "0110000101110100" when "1010111001",
   "0110000110010000" when "1010111010",
   "0110000110101011" when "1010111011",
   "0110000111000111" when "1010111100",
   "0110000111100011" when "1010111101",
   "0110000111111111" when "1010111110",
   "0110001000011010" when "1010111111",
   "0110001000110110" when "1011000000",
   "0110001001010010" when "1011000001",
   "0110001001101101" when "1011000010",
   "0110001010001001" when "1011000011",
   "0110001010100100" when "1011000100",
   "0110001011000000" when "1011000101",
   "0110001011011011" when "1011000110",
   "0110001011110111" when "1011000111",
   "0110001100010010" when "1011001000",
   "0110001100101110" when "1011001001",
   "0110001101001001" when "1011001010",
   "0110001101100101" when "1011001011",
   "0110001110000000" when "1011001100",
   "0110001110011011" when "1011001101",
   "0110001110110111" when "1011001110",
   "0110001111010010" when "1011001111",
   "0110001111101101" when "1011010000",
   "0110010000001000" when "1011010001",
   "0110010000100100" when "1011010010",
   "0110010000111111" when "1011010011",
   "0110010001011010" when "1011010100",
   "0110010001110101" when "1011010101",
   "0110010010010000" when "1011010110",
   "0110010010101011" when "1011010111",
   "0110010011000110" when "1011011000",
   "0110010011100001" when "1011011001",
   "0110010011111100" when "1011011010",
   "0110010100010111" when "1011011011",
   "0110010100110010" when "1011011100",
   "0110010101001101" when "1011011101",
   "0110010101101000" when "1011011110",
   "0110010110000011" when "1011011111",
   "0110010110011110" when "1011100000",
   "0110010110111001" when "1011100001",
   "0110010111010100" when "1011100010",
   "0110010111101110" when "1011100011",
   "0110011000001001" when "1011100100",
   "0110011000100100" when "1011100101",
   "0110011000111111" when "1011100110",
   "0110011001011001" when "1011100111",
   "0110011001110100" when "1011101000",
   "0110011010001111" when "1011101001",
   "0110011010101001" when "1011101010",
   "0110011011000100" when "1011101011",
   "0110011011011110" when "1011101100",
   "0110011011111001" when "1011101101",
   "0110011100010100" when "1011101110",
   "0110011100101110" when "1011101111",
   "0110011101001001" when "1011110000",
   "0110011101100011" when "1011110001",
   "0110011101111101" when "1011110010",
   "0110011110011000" when "1011110011",
   "0110011110110010" when "1011110100",
   "0110011111001100" when "1011110101",
   "0110011111100111" when "1011110110",
   "0110100000000001" when "1011110111",
   "0110100000011011" when "1011111000",
   "0110100000110110" when "1011111001",
   "0110100001010000" when "1011111010",
   "0110100001101010" when "1011111011",
   "0110100010000100" when "1011111100",
   "0110100010011110" when "1011111101",
   "0110100010111000" when "1011111110",
   "0110100011010011" when "1011111111",
   "0110100011101101" when "1100000000",
   "0110100100000111" when "1100000001",
   "0110100100100001" when "1100000010",
   "0110100100111011" when "1100000011",
   "0110100101010101" when "1100000100",
   "0110100101101111" when "1100000101",
   "0110100110001001" when "1100000110",
   "0110100110100011" when "1100000111",
   "0110100110111100" when "1100001000",
   "0110100111010110" when "1100001001",
   "0110100111110000" when "1100001010",
   "0110101000001010" when "1100001011",
   "0110101000100100" when "1100001100",
   "0110101000111101" when "1100001101",
   "0110101001010111" when "1100001110",
   "0110101001110001" when "1100001111",
   "0110101010001011" when "1100010000",
   "0110101010100100" when "1100010001",
   "0110101010111110" when "1100010010",
   "0110101011010111" when "1100010011",
   "0110101011110001" when "1100010100",
   "0110101100001011" when "1100010101",
   "0110101100100100" when "1100010110",
   "0110101100111110" when "1100010111",
   "0110101101010111" when "1100011000",
   "0110101101110001" when "1100011001",
   "0110101110001010" when "1100011010",
   "0110101110100100" when "1100011011",
   "0110101110111101" when "1100011100",
   "0110101111010110" when "1100011101",
   "0110101111110000" when "1100011110",
   "0110110000001001" when "1100011111",
   "0110110000100010" when "1100100000",
   "0110110000111100" when "1100100001",
   "0110110001010101" when "1100100010",
   "0110110001101110" when "1100100011",
   "0110110010000111" when "1100100100",
   "0110110010100000" when "1100100101",
   "0110110010111010" when "1100100110",
   "0110110011010011" when "1100100111",
   "0110110011101100" when "1100101000",
   "0110110100000101" when "1100101001",
   "0110110100011110" when "1100101010",
   "0110110100110111" when "1100101011",
   "0110110101010000" when "1100101100",
   "0110110101101001" when "1100101101",
   "0110110110000010" when "1100101110",
   "0110110110011011" when "1100101111",
   "0110110110110100" when "1100110000",
   "0110110111001101" when "1100110001",
   "0110110111100110" when "1100110010",
   "0110110111111110" when "1100110011",
   "0110111000010111" when "1100110100",
   "0110111000110000" when "1100110101",
   "0110111001001001" when "1100110110",
   "0110111001100010" when "1100110111",
   "0110111001111010" when "1100111000",
   "0110111010010011" when "1100111001",
   "0110111010101100" when "1100111010",
   "0110111011000100" when "1100111011",
   "0110111011011101" when "1100111100",
   "0110111011110110" when "1100111101",
   "0110111100001110" when "1100111110",
   "0110111100100111" when "1100111111",
   "0110111100111111" when "1101000000",
   "0110111101011000" when "1101000001",
   "0110111101110000" when "1101000010",
   "0110111110001001" when "1101000011",
   "0110111110100001" when "1101000100",
   "0110111110111010" when "1101000101",
   "0110111111010010" when "1101000110",
   "0110111111101010" when "1101000111",
   "0111000000000011" when "1101001000",
   "0111000000011011" when "1101001001",
   "0111000000110011" when "1101001010",
   "0111000001001100" when "1101001011",
   "0111000001100100" when "1101001100",
   "0111000001111100" when "1101001101",
   "0111000010010100" when "1101001110",
   "0111000010101101" when "1101001111",
   "0111000011000101" when "1101010000",
   "0111000011011101" when "1101010001",
   "0111000011110101" when "1101010010",
   "0111000100001101" when "1101010011",
   "0111000100100101" when "1101010100",
   "0111000100111101" when "1101010101",
   "0111000101010101" when "1101010110",
   "0111000101101101" when "1101010111",
   "0111000110000101" when "1101011000",
   "0111000110011101" when "1101011001",
   "0111000110110101" when "1101011010",
   "0111000111001101" when "1101011011",
   "0111000111100101" when "1101011100",
   "0111000111111101" when "1101011101",
   "0111001000010101" when "1101011110",
   "0111001000101101" when "1101011111",
   "0111001001000100" when "1101100000",
   "0111001001011100" when "1101100001",
   "0111001001110100" when "1101100010",
   "0111001010001100" when "1101100011",
   "0111001010100011" when "1101100100",
   "0111001010111011" when "1101100101",
   "0111001011010011" when "1101100110",
   "0111001011101010" when "1101100111",
   "0111001100000010" when "1101101000",
   "0111001100011010" when "1101101001",
   "0111001100110001" when "1101101010",
   "0111001101001001" when "1101101011",
   "0111001101100000" when "1101101100",
   "0111001101111000" when "1101101101",
   "0111001110001111" when "1101101110",
   "0111001110100111" when "1101101111",
   "0111001110111110" when "1101110000",
   "0111001111010110" when "1101110001",
   "0111001111101101" when "1101110010",
   "0111010000000100" when "1101110011",
   "0111010000011100" when "1101110100",
   "0111010000110011" when "1101110101",
   "0111010001001010" when "1101110110",
   "0111010001100010" when "1101110111",
   "0111010001111001" when "1101111000",
   "0111010010010000" when "1101111001",
   "0111010010100111" when "1101111010",
   "0111010010111110" when "1101111011",
   "0111010011010110" when "1101111100",
   "0111010011101101" when "1101111101",
   "0111010100000100" when "1101111110",
   "0111010100011011" when "1101111111",
   "0111010100110010" when "1110000000",
   "0111010101001001" when "1110000001",
   "0111010101100000" when "1110000010",
   "0111010101110111" when "1110000011",
   "0111010110001110" when "1110000100",
   "0111010110100101" when "1110000101",
   "0111010110111100" when "1110000110",
   "0111010111010011" when "1110000111",
   "0111010111101010" when "1110001000",
   "0111011000000001" when "1110001001",
   "0111011000011000" when "1110001010",
   "0111011000101110" when "1110001011",
   "0111011001000101" when "1110001100",
   "0111011001011100" when "1110001101",
   "0111011001110011" when "1110001110",
   "0111011010001010" when "1110001111",
   "0111011010100000" when "1110010000",
   "0111011010110111" when "1110010001",
   "0111011011001110" when "1110010010",
   "0111011011100100" when "1110010011",
   "0111011011111011" when "1110010100",
   "0111011100010010" when "1110010101",
   "0111011100101000" when "1110010110",
   "0111011100111111" when "1110010111",
   "0111011101010101" when "1110011000",
   "0111011101101100" when "1110011001",
   "0111011110000010" when "1110011010",
   "0111011110011001" when "1110011011",
   "0111011110101111" when "1110011100",
   "0111011111000110" when "1110011101",
   "0111011111011100" when "1110011110",
   "0111011111110010" when "1110011111",
   "0111100000001001" when "1110100000",
   "0111100000011111" when "1110100001",
   "0111100000110101" when "1110100010",
   "0111100001001100" when "1110100011",
   "0111100001100010" when "1110100100",
   "0111100001111000" when "1110100101",
   "0111100010001111" when "1110100110",
   "0111100010100101" when "1110100111",
   "0111100010111011" when "1110101000",
   "0111100011010001" when "1110101001",
   "0111100011100111" when "1110101010",
   "0111100011111101" when "1110101011",
   "0111100100010100" when "1110101100",
   "0111100100101010" when "1110101101",
   "0111100101000000" when "1110101110",
   "0111100101010110" when "1110101111",
   "0111100101101100" when "1110110000",
   "0111100110000010" when "1110110001",
   "0111100110011000" when "1110110010",
   "0111100110101110" when "1110110011",
   "0111100111000100" when "1110110100",
   "0111100111011010" when "1110110101",
   "0111100111101111" when "1110110110",
   "0111101000000101" when "1110110111",
   "0111101000011011" when "1110111000",
   "0111101000110001" when "1110111001",
   "0111101001000111" when "1110111010",
   "0111101001011101" when "1110111011",
   "0111101001110010" when "1110111100",
   "0111101010001000" when "1110111101",
   "0111101010011110" when "1110111110",
   "0111101010110100" when "1110111111",
   "0111101011001001" when "1111000000",
   "0111101011011111" when "1111000001",
   "0111101011110101" when "1111000010",
   "0111101100001010" when "1111000011",
   "0111101100100000" when "1111000100",
   "0111101100110101" when "1111000101",
   "0111101101001011" when "1111000110",
   "0111101101100000" when "1111000111",
   "0111101101110110" when "1111001000",
   "0111101110001011" when "1111001001",
   "0111101110100001" when "1111001010",
   "0111101110110110" when "1111001011",
   "0111101111001100" when "1111001100",
   "0111101111100001" when "1111001101",
   "0111101111110111" when "1111001110",
   "0111110000001100" when "1111001111",
   "0111110000100001" when "1111010000",
   "0111110000110111" when "1111010001",
   "0111110001001100" when "1111010010",
   "0111110001100001" when "1111010011",
   "0111110001110111" when "1111010100",
   "0111110010001100" when "1111010101",
   "0111110010100001" when "1111010110",
   "0111110010110110" when "1111010111",
   "0111110011001011" when "1111011000",
   "0111110011100001" when "1111011001",
   "0111110011110110" when "1111011010",
   "0111110100001011" when "1111011011",
   "0111110100100000" when "1111011100",
   "0111110100110101" when "1111011101",
   "0111110101001010" when "1111011110",
   "0111110101011111" when "1111011111",
   "0111110101110100" when "1111100000",
   "0111110110001001" when "1111100001",
   "0111110110011110" when "1111100010",
   "0111110110110011" when "1111100011",
   "0111110111001000" when "1111100100",
   "0111110111011101" when "1111100101",
   "0111110111110010" when "1111100110",
   "0111111000000111" when "1111100111",
   "0111111000011100" when "1111101000",
   "0111111000110000" when "1111101001",
   "0111111001000101" when "1111101010",
   "0111111001011010" when "1111101011",
   "0111111001101111" when "1111101100",
   "0111111010000100" when "1111101101",
   "0111111010011000" when "1111101110",
   "0111111010101101" when "1111101111",
   "0111111011000010" when "1111110000",
   "0111111011010110" when "1111110001",
   "0111111011101011" when "1111110010",
   "0111111100000000" when "1111110011",
   "0111111100010100" when "1111110100",
   "0111111100101001" when "1111110101",
   "0111111100111101" when "1111110110",
   "0111111101010010" when "1111110111",
   "0111111101100110" when "1111111000",
   "0111111101111011" when "1111111001",
   "0111111110001111" when "1111111010",
   "0111111110100100" when "1111111011",
   "0111111110111000" when "1111111100",
   "0111111111001101" when "1111111101",
   "0111111111100001" when "1111111110",
   "0111111111110110" when "1111111111",
   "----------------" when others;
    Y <= TableOut_d1;
end architecture;

--------------------------------------------------------------------------------
--                        GenericTable_10_6_F400_uid33
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity GenericTable_10_6_F400_uid33 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(9 downto 0);
          Y : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericTable_10_6_F400_uid33 is
signal TableOut :  std_logic_vector(5 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
  with X select TableOut <= 
   "101100" when "0000000000",
   "101101" when "0000000001",
   "101101" when "0000000010",
   "101110" when "0000000011",
   "101110" when "0000000100",
   "101111" when "0000000101",
   "110000" when "0000000110",
   "110000" when "0000000111",
   "110001" when "0000001000",
   "110010" when "0000001001",
   "110010" when "0000001010",
   "110011" when "0000001011",
   "110100" when "0000001100",
   "110100" when "0000001101",
   "110101" when "0000001110",
   "110101" when "0000001111",
   "110110" when "0000010000",
   "110111" when "0000010001",
   "110111" when "0000010010",
   "111000" when "0000010011",
   "111001" when "0000010100",
   "111001" when "0000010101",
   "111010" when "0000010110",
   "111011" when "0000010111",
   "111011" when "0000011000",
   "111100" when "0000011001",
   "111100" when "0000011010",
   "111101" when "0000011011",
   "111110" when "0000011100",
   "111110" when "0000011101",
   "111111" when "0000011110",
   "111111" when "0000011111",
   "101100" when "0000100000",
   "101101" when "0000100001",
   "101101" when "0000100010",
   "101110" when "0000100011",
   "101111" when "0000100100",
   "101111" when "0000100101",
   "110000" when "0000100110",
   "110000" when "0000100111",
   "110001" when "0000101000",
   "110010" when "0000101001",
   "110010" when "0000101010",
   "110011" when "0000101011",
   "110100" when "0000101100",
   "110100" when "0000101101",
   "110101" when "0000101110",
   "110110" when "0000101111",
   "110110" when "0000110000",
   "110111" when "0000110001",
   "110111" when "0000110010",
   "111000" when "0000110011",
   "111001" when "0000110100",
   "111001" when "0000110101",
   "111010" when "0000110110",
   "111011" when "0000110111",
   "111011" when "0000111000",
   "111100" when "0000111001",
   "111101" when "0000111010",
   "111101" when "0000111011",
   "111110" when "0000111100",
   "111110" when "0000111101",
   "111111" when "0000111110",
   "111111" when "0000111111",
   "101100" when "0001000000",
   "101101" when "0001000001",
   "101101" when "0001000010",
   "101110" when "0001000011",
   "101111" when "0001000100",
   "101111" when "0001000101",
   "110000" when "0001000110",
   "110000" when "0001000111",
   "110001" when "0001001000",
   "110010" when "0001001001",
   "110010" when "0001001010",
   "110011" when "0001001011",
   "110100" when "0001001100",
   "110100" when "0001001101",
   "110101" when "0001001110",
   "110110" when "0001001111",
   "110110" when "0001010000",
   "110111" when "0001010001",
   "110111" when "0001010010",
   "111000" when "0001010011",
   "111001" when "0001010100",
   "111001" when "0001010101",
   "111010" when "0001010110",
   "111011" when "0001010111",
   "111011" when "0001011000",
   "111100" when "0001011001",
   "111101" when "0001011010",
   "111101" when "0001011011",
   "111110" when "0001011100",
   "111110" when "0001011101",
   "111111" when "0001011110",
   "111111" when "0001011111",
   "101100" when "0001100000",
   "101101" when "0001100001",
   "101101" when "0001100010",
   "101110" when "0001100011",
   "101111" when "0001100100",
   "101111" when "0001100101",
   "110000" when "0001100110",
   "110001" when "0001100111",
   "110001" when "0001101000",
   "110010" when "0001101001",
   "110010" when "0001101010",
   "110011" when "0001101011",
   "110100" when "0001101100",
   "110100" when "0001101101",
   "110101" when "0001101110",
   "110110" when "0001101111",
   "110110" when "0001110000",
   "110111" when "0001110001",
   "111000" when "0001110010",
   "111000" when "0001110011",
   "111001" when "0001110100",
   "111001" when "0001110101",
   "111010" when "0001110110",
   "111011" when "0001110111",
   "111011" when "0001111000",
   "111100" when "0001111001",
   "111101" when "0001111010",
   "111101" when "0001111011",
   "111110" when "0001111100",
   "111110" when "0001111101",
   "111111" when "0001111110",
   "111111" when "0001111111",
   "101100" when "0010000000",
   "101101" when "0010000001",
   "101110" when "0010000010",
   "101110" when "0010000011",
   "101111" when "0010000100",
   "101111" when "0010000101",
   "110000" when "0010000110",
   "110001" when "0010000111",
   "110001" when "0010001000",
   "110010" when "0010001001",
   "110011" when "0010001010",
   "110011" when "0010001011",
   "110100" when "0010001100",
   "110100" when "0010001101",
   "110101" when "0010001110",
   "110110" when "0010001111",
   "110110" when "0010010000",
   "110111" when "0010010001",
   "111000" when "0010010010",
   "111000" when "0010010011",
   "111001" when "0010010100",
   "111001" when "0010010101",
   "111010" when "0010010110",
   "111011" when "0010010111",
   "111011" when "0010011000",
   "111100" when "0010011001",
   "111101" when "0010011010",
   "111101" when "0010011011",
   "111110" when "0010011100",
   "111110" when "0010011101",
   "111111" when "0010011110",
   "111111" when "0010011111",
   "101101" when "0010100000",
   "101101" when "0010100001",
   "101110" when "0010100010",
   "101110" when "0010100011",
   "101111" when "0010100100",
   "110000" when "0010100101",
   "110000" when "0010100110",
   "110001" when "0010100111",
   "110001" when "0010101000",
   "110010" when "0010101001",
   "110011" when "0010101010",
   "110011" when "0010101011",
   "110100" when "0010101100",
   "110101" when "0010101101",
   "110101" when "0010101110",
   "110110" when "0010101111",
   "110110" when "0010110000",
   "110111" when "0010110001",
   "111000" when "0010110010",
   "111000" when "0010110011",
   "111001" when "0010110100",
   "111010" when "0010110101",
   "111010" when "0010110110",
   "111011" when "0010110111",
   "111011" when "0010111000",
   "111100" when "0010111001",
   "111101" when "0010111010",
   "111101" when "0010111011",
   "111110" when "0010111100",
   "111110" when "0010111101",
   "111111" when "0010111110",
   "111111" when "0010111111",
   "101101" when "0011000000",
   "101101" when "0011000001",
   "101110" when "0011000010",
   "101111" when "0011000011",
   "101111" when "0011000100",
   "110000" when "0011000101",
   "110000" when "0011000110",
   "110001" when "0011000111",
   "110010" when "0011001000",
   "110010" when "0011001001",
   "110011" when "0011001010",
   "110011" when "0011001011",
   "110100" when "0011001100",
   "110101" when "0011001101",
   "110101" when "0011001110",
   "110110" when "0011001111",
   "110111" when "0011010000",
   "110111" when "0011010001",
   "111000" when "0011010010",
   "111000" when "0011010011",
   "111001" when "0011010100",
   "111010" when "0011010101",
   "111010" when "0011010110",
   "111011" when "0011010111",
   "111011" when "0011011000",
   "111100" when "0011011001",
   "111101" when "0011011010",
   "111101" when "0011011011",
   "111110" when "0011011100",
   "111110" when "0011011101",
   "111111" when "0011011110",
   "111111" when "0011011111",
   "101101" when "0011100000",
   "101110" when "0011100001",
   "101110" when "0011100010",
   "101111" when "0011100011",
   "101111" when "0011100100",
   "110000" when "0011100101",
   "110001" when "0011100110",
   "110001" when "0011100111",
   "110010" when "0011101000",
   "110010" when "0011101001",
   "110011" when "0011101010",
   "110100" when "0011101011",
   "110100" when "0011101100",
   "110101" when "0011101101",
   "110101" when "0011101110",
   "110110" when "0011101111",
   "110111" when "0011110000",
   "110111" when "0011110001",
   "111000" when "0011110010",
   "111000" when "0011110011",
   "111001" when "0011110100",
   "111010" when "0011110101",
   "111010" when "0011110110",
   "111011" when "0011110111",
   "111011" when "0011111000",
   "111100" when "0011111001",
   "111101" when "0011111010",
   "111101" when "0011111011",
   "111110" when "0011111100",
   "111110" when "0011111101",
   "111111" when "0011111110",
   "111111" when "0011111111",
   "101101" when "0100000000",
   "101110" when "0100000001",
   "101110" when "0100000010",
   "101111" when "0100000011",
   "110000" when "0100000100",
   "110000" when "0100000101",
   "110001" when "0100000110",
   "110001" when "0100000111",
   "110010" when "0100001000",
   "110011" when "0100001001",
   "110011" when "0100001010",
   "110100" when "0100001011",
   "110100" when "0100001100",
   "110101" when "0100001101",
   "110110" when "0100001110",
   "110110" when "0100001111",
   "110111" when "0100010000",
   "110111" when "0100010001",
   "111000" when "0100010010",
   "111001" when "0100010011",
   "111001" when "0100010100",
   "111010" when "0100010101",
   "111010" when "0100010110",
   "111011" when "0100010111",
   "111100" when "0100011000",
   "111100" when "0100011001",
   "111101" when "0100011010",
   "111101" when "0100011011",
   "111110" when "0100011100",
   "111111" when "0100011101",
   "111111" when "0100011110",
   "111111" when "0100011111",
   "101110" when "0100100000",
   "101110" when "0100100001",
   "101111" when "0100100010",
   "101111" when "0100100011",
   "110000" when "0100100100",
   "110000" when "0100100101",
   "110001" when "0100100110",
   "110010" when "0100100111",
   "110010" when "0100101000",
   "110011" when "0100101001",
   "110011" when "0100101010",
   "110100" when "0100101011",
   "110101" when "0100101100",
   "110101" when "0100101101",
   "110110" when "0100101110",
   "110110" when "0100101111",
   "110111" when "0100110000",
   "111000" when "0100110001",
   "111000" when "0100110010",
   "111001" when "0100110011",
   "111001" when "0100110100",
   "111010" when "0100110101",
   "111010" when "0100110110",
   "111011" when "0100110111",
   "111100" when "0100111000",
   "111100" when "0100111001",
   "111101" when "0100111010",
   "111101" when "0100111011",
   "111110" when "0100111100",
   "111111" when "0100111101",
   "111111" when "0100111110",
   "111111" when "0100111111",
   "101110" when "0101000000",
   "101110" when "0101000001",
   "101111" when "0101000010",
   "110000" when "0101000011",
   "110000" when "0101000100",
   "110001" when "0101000101",
   "110001" when "0101000110",
   "110010" when "0101000111",
   "110010" when "0101001000",
   "110011" when "0101001001",
   "110100" when "0101001010",
   "110100" when "0101001011",
   "110101" when "0101001100",
   "110101" when "0101001101",
   "110110" when "0101001110",
   "110111" when "0101001111",
   "110111" when "0101010000",
   "111000" when "0101010001",
   "111000" when "0101010010",
   "111001" when "0101010011",
   "111001" when "0101010100",
   "111010" when "0101010101",
   "111011" when "0101010110",
   "111011" when "0101010111",
   "111100" when "0101011000",
   "111100" when "0101011001",
   "111101" when "0101011010",
   "111101" when "0101011011",
   "111110" when "0101011100",
   "111111" when "0101011101",
   "111111" when "0101011110",
   "111111" when "0101011111",
   "101110" when "0101100000",
   "101111" when "0101100001",
   "101111" when "0101100010",
   "110000" when "0101100011",
   "110000" when "0101100100",
   "110001" when "0101100101",
   "110010" when "0101100110",
   "110010" when "0101100111",
   "110011" when "0101101000",
   "110011" when "0101101001",
   "110100" when "0101101010",
   "110100" when "0101101011",
   "110101" when "0101101100",
   "110110" when "0101101101",
   "110110" when "0101101110",
   "110111" when "0101101111",
   "110111" when "0101110000",
   "111000" when "0101110001",
   "111000" when "0101110010",
   "111001" when "0101110011",
   "111010" when "0101110100",
   "111010" when "0101110101",
   "111011" when "0101110110",
   "111011" when "0101110111",
   "111100" when "0101111000",
   "111100" when "0101111001",
   "111101" when "0101111010",
   "111101" when "0101111011",
   "111110" when "0101111100",
   "111111" when "0101111101",
   "111111" when "0101111110",
   "111111" when "0101111111",
   "101111" when "0110000000",
   "101111" when "0110000001",
   "110000" when "0110000010",
   "110000" when "0110000011",
   "110001" when "0110000100",
   "110001" when "0110000101",
   "110010" when "0110000110",
   "110010" when "0110000111",
   "110011" when "0110001000",
   "110100" when "0110001001",
   "110100" when "0110001010",
   "110101" when "0110001011",
   "110101" when "0110001100",
   "110110" when "0110001101",
   "110110" when "0110001110",
   "110111" when "0110001111",
   "110111" when "0110010000",
   "111000" when "0110010001",
   "111001" when "0110010010",
   "111001" when "0110010011",
   "111010" when "0110010100",
   "111010" when "0110010101",
   "111011" when "0110010110",
   "111011" when "0110010111",
   "111100" when "0110011000",
   "111100" when "0110011001",
   "111101" when "0110011010",
   "111110" when "0110011011",
   "111110" when "0110011100",
   "111111" when "0110011101",
   "111111" when "0110011110",
   "111111" when "0110011111",
   "101111" when "0110100000",
   "110000" when "0110100001",
   "110000" when "0110100010",
   "110001" when "0110100011",
   "110001" when "0110100100",
   "110010" when "0110100101",
   "110010" when "0110100110",
   "110011" when "0110100111",
   "110011" when "0110101000",
   "110100" when "0110101001",
   "110100" when "0110101010",
   "110101" when "0110101011",
   "110101" when "0110101100",
   "110110" when "0110101101",
   "110111" when "0110101110",
   "110111" when "0110101111",
   "111000" when "0110110000",
   "111000" when "0110110001",
   "111001" when "0110110010",
   "111001" when "0110110011",
   "111010" when "0110110100",
   "111010" when "0110110101",
   "111011" when "0110110110",
   "111011" when "0110110111",
   "111100" when "0110111000",
   "111100" when "0110111001",
   "111101" when "0110111010",
   "111110" when "0110111011",
   "111110" when "0110111100",
   "111111" when "0110111101",
   "111111" when "0110111110",
   "111111" when "0110111111",
   "101111" when "0111000000",
   "110000" when "0111000001",
   "110000" when "0111000010",
   "110001" when "0111000011",
   "110001" when "0111000100",
   "110010" when "0111000101",
   "110011" when "0111000110",
   "110011" when "0111000111",
   "110100" when "0111001000",
   "110100" when "0111001001",
   "110101" when "0111001010",
   "110101" when "0111001011",
   "110110" when "0111001100",
   "110110" when "0111001101",
   "110111" when "0111001110",
   "110111" when "0111001111",
   "111000" when "0111010000",
   "111000" when "0111010001",
   "111001" when "0111010010",
   "111001" when "0111010011",
   "111010" when "0111010100",
   "111010" when "0111010101",
   "111011" when "0111010110",
   "111100" when "0111010111",
   "111100" when "0111011000",
   "111101" when "0111011001",
   "111101" when "0111011010",
   "111110" when "0111011011",
   "111110" when "0111011100",
   "111111" when "0111011101",
   "111111" when "0111011110",
   "111111" when "0111011111",
   "110000" when "0111100000",
   "110000" when "0111100001",
   "110001" when "0111100010",
   "110001" when "0111100011",
   "110010" when "0111100100",
   "110010" when "0111100101",
   "110011" when "0111100110",
   "110011" when "0111100111",
   "110100" when "0111101000",
   "110100" when "0111101001",
   "110101" when "0111101010",
   "110101" when "0111101011",
   "110110" when "0111101100",
   "110110" when "0111101101",
   "110111" when "0111101110",
   "110111" when "0111101111",
   "111000" when "0111110000",
   "111001" when "0111110001",
   "111001" when "0111110010",
   "111010" when "0111110011",
   "111010" when "0111110100",
   "111011" when "0111110101",
   "111011" when "0111110110",
   "111100" when "0111110111",
   "111100" when "0111111000",
   "111101" when "0111111001",
   "111101" when "0111111010",
   "111110" when "0111111011",
   "111110" when "0111111100",
   "111111" when "0111111101",
   "111111" when "0111111110",
   "111111" when "0111111111",
   "110000" when "1000000000",
   "110001" when "1000000001",
   "110001" when "1000000010",
   "110010" when "1000000011",
   "110010" when "1000000100",
   "110011" when "1000000101",
   "110011" when "1000000110",
   "110100" when "1000000111",
   "110100" when "1000001000",
   "110101" when "1000001001",
   "110101" when "1000001010",
   "110110" when "1000001011",
   "110110" when "1000001100",
   "110111" when "1000001101",
   "110111" when "1000001110",
   "111000" when "1000001111",
   "111000" when "1000010000",
   "111001" when "1000010001",
   "111001" when "1000010010",
   "111010" when "1000010011",
   "111010" when "1000010100",
   "111011" when "1000010101",
   "111011" when "1000010110",
   "111100" when "1000010111",
   "111100" when "1000011000",
   "111101" when "1000011001",
   "111101" when "1000011010",
   "111110" when "1000011011",
   "111110" when "1000011100",
   "111111" when "1000011101",
   "111111" when "1000011110",
   "111111" when "1000011111",
   "110001" when "1000100000",
   "110001" when "1000100001",
   "110010" when "1000100010",
   "110010" when "1000100011",
   "110011" when "1000100100",
   "110011" when "1000100101",
   "110100" when "1000100110",
   "110100" when "1000100111",
   "110100" when "1000101000",
   "110101" when "1000101001",
   "110101" when "1000101010",
   "110110" when "1000101011",
   "110110" when "1000101100",
   "110111" when "1000101101",
   "110111" when "1000101110",
   "111000" when "1000101111",
   "111000" when "1000110000",
   "111001" when "1000110001",
   "111001" when "1000110010",
   "111010" when "1000110011",
   "111010" when "1000110100",
   "111011" when "1000110101",
   "111011" when "1000110110",
   "111100" when "1000110111",
   "111100" when "1000111000",
   "111101" when "1000111001",
   "111101" when "1000111010",
   "111110" when "1000111011",
   "111110" when "1000111100",
   "111111" when "1000111101",
   "111111" when "1000111110",
   "111111" when "1000111111",
   "110001" when "1001000000",
   "110001" when "1001000001",
   "110010" when "1001000010",
   "110010" when "1001000011",
   "110011" when "1001000100",
   "110011" when "1001000101",
   "110100" when "1001000110",
   "110100" when "1001000111",
   "110101" when "1001001000",
   "110101" when "1001001001",
   "110110" when "1001001010",
   "110110" when "1001001011",
   "110111" when "1001001100",
   "110111" when "1001001101",
   "111000" when "1001001110",
   "111000" when "1001001111",
   "111001" when "1001010000",
   "111001" when "1001010001",
   "111010" when "1001010010",
   "111010" when "1001010011",
   "111011" when "1001010100",
   "111011" when "1001010101",
   "111011" when "1001010110",
   "111100" when "1001010111",
   "111100" when "1001011000",
   "111101" when "1001011001",
   "111101" when "1001011010",
   "111110" when "1001011011",
   "111110" when "1001011100",
   "111111" when "1001011101",
   "111111" when "1001011110",
   "111111" when "1001011111",
   "110001" when "1001100000",
   "110010" when "1001100001",
   "110010" when "1001100010",
   "110011" when "1001100011",
   "110011" when "1001100100",
   "110100" when "1001100101",
   "110100" when "1001100110",
   "110101" when "1001100111",
   "110101" when "1001101000",
   "110110" when "1001101001",
   "110110" when "1001101010",
   "110110" when "1001101011",
   "110111" when "1001101100",
   "110111" when "1001101101",
   "111000" when "1001101110",
   "111000" when "1001101111",
   "111001" when "1001110000",
   "111001" when "1001110001",
   "111010" when "1001110010",
   "111010" when "1001110011",
   "111011" when "1001110100",
   "111011" when "1001110101",
   "111100" when "1001110110",
   "111100" when "1001110111",
   "111101" when "1001111000",
   "111101" when "1001111001",
   "111101" when "1001111010",
   "111110" when "1001111011",
   "111110" when "1001111100",
   "111111" when "1001111101",
   "111111" when "1001111110",
   "111111" when "1001111111",
   "110010" when "1010000000",
   "110010" when "1010000001",
   "110011" when "1010000010",
   "110011" when "1010000011",
   "110100" when "1010000100",
   "110100" when "1010000101",
   "110100" when "1010000110",
   "110101" when "1010000111",
   "110101" when "1010001000",
   "110110" when "1010001001",
   "110110" when "1010001010",
   "110111" when "1010001011",
   "110111" when "1010001100",
   "111000" when "1010001101",
   "111000" when "1010001110",
   "111001" when "1010001111",
   "111001" when "1010010000",
   "111001" when "1010010001",
   "111010" when "1010010010",
   "111010" when "1010010011",
   "111011" when "1010010100",
   "111011" when "1010010101",
   "111100" when "1010010110",
   "111100" when "1010010111",
   "111101" when "1010011000",
   "111101" when "1010011001",
   "111110" when "1010011010",
   "111110" when "1010011011",
   "111110" when "1010011100",
   "111111" when "1010011101",
   "111111" when "1010011110",
   "111111" when "1010011111",
   "110010" when "1010100000",
   "110011" when "1010100001",
   "110011" when "1010100010",
   "110011" when "1010100011",
   "110100" when "1010100100",
   "110100" when "1010100101",
   "110101" when "1010100110",
   "110101" when "1010100111",
   "110110" when "1010101000",
   "110110" when "1010101001",
   "110111" when "1010101010",
   "110111" when "1010101011",
   "110111" when "1010101100",
   "111000" when "1010101101",
   "111000" when "1010101110",
   "111001" when "1010101111",
   "111001" when "1010110000",
   "111010" when "1010110001",
   "111010" when "1010110010",
   "111011" when "1010110011",
   "111011" when "1010110100",
   "111011" when "1010110101",
   "111100" when "1010110110",
   "111100" when "1010110111",
   "111101" when "1010111000",
   "111101" when "1010111001",
   "111110" when "1010111010",
   "111110" when "1010111011",
   "111110" when "1010111100",
   "111111" when "1010111101",
   "111111" when "1010111110",
   "111111" when "1010111111",
   "110011" when "1011000000",
   "110011" when "1011000001",
   "110011" when "1011000010",
   "110100" when "1011000011",
   "110100" when "1011000100",
   "110101" when "1011000101",
   "110101" when "1011000110",
   "110110" when "1011000111",
   "110110" when "1011001000",
   "110110" when "1011001001",
   "110111" when "1011001010",
   "110111" when "1011001011",
   "111000" when "1011001100",
   "111000" when "1011001101",
   "111001" when "1011001110",
   "111001" when "1011001111",
   "111001" when "1011010000",
   "111010" when "1011010001",
   "111010" when "1011010010",
   "111011" when "1011010011",
   "111011" when "1011010100",
   "111100" when "1011010101",
   "111100" when "1011010110",
   "111100" when "1011010111",
   "111101" when "1011011000",
   "111101" when "1011011001",
   "111110" when "1011011010",
   "111110" when "1011011011",
   "111111" when "1011011100",
   "111111" when "1011011101",
   "111111" when "1011011110",
   "111111" when "1011011111",
   "110011" when "1011100000",
   "110011" when "1011100001",
   "110100" when "1011100010",
   "110100" when "1011100011",
   "110101" when "1011100100",
   "110101" when "1011100101",
   "110101" when "1011100110",
   "110110" when "1011100111",
   "110110" when "1011101000",
   "110111" when "1011101001",
   "110111" when "1011101010",
   "111000" when "1011101011",
   "111000" when "1011101100",
   "111000" when "1011101101",
   "111001" when "1011101110",
   "111001" when "1011101111",
   "111010" when "1011110000",
   "111010" when "1011110001",
   "111010" when "1011110010",
   "111011" when "1011110011",
   "111011" when "1011110100",
   "111100" when "1011110101",
   "111100" when "1011110110",
   "111100" when "1011110111",
   "111101" when "1011111000",
   "111101" when "1011111001",
   "111110" when "1011111010",
   "111110" when "1011111011",
   "111111" when "1011111100",
   "111111" when "1011111101",
   "111111" when "1011111110",
   "111111" when "1011111111",
   "110011" when "1100000000",
   "110100" when "1100000001",
   "110100" when "1100000010",
   "110101" when "1100000011",
   "110101" when "1100000100",
   "110101" when "1100000101",
   "110110" when "1100000110",
   "110110" when "1100000111",
   "110111" when "1100001000",
   "110111" when "1100001001",
   "110111" when "1100001010",
   "111000" when "1100001011",
   "111000" when "1100001100",
   "111001" when "1100001101",
   "111001" when "1100001110",
   "111001" when "1100001111",
   "111010" when "1100010000",
   "111010" when "1100010001",
   "111011" when "1100010010",
   "111011" when "1100010011",
   "111011" when "1100010100",
   "111100" when "1100010101",
   "111100" when "1100010110",
   "111101" when "1100010111",
   "111101" when "1100011000",
   "111101" when "1100011001",
   "111110" when "1100011010",
   "111110" when "1100011011",
   "111111" when "1100011100",
   "111111" when "1100011101",
   "111111" when "1100011110",
   "111111" when "1100011111",
   "110100" when "1100100000",
   "110100" when "1100100001",
   "110101" when "1100100010",
   "110101" when "1100100011",
   "110101" when "1100100100",
   "110110" when "1100100101",
   "110110" when "1100100110",
   "110110" when "1100100111",
   "110111" when "1100101000",
   "110111" when "1100101001",
   "111000" when "1100101010",
   "111000" when "1100101011",
   "111000" when "1100101100",
   "111001" when "1100101101",
   "111001" when "1100101110",
   "111010" when "1100101111",
   "111010" when "1100110000",
   "111010" when "1100110001",
   "111011" when "1100110010",
   "111011" when "1100110011",
   "111100" when "1100110100",
   "111100" when "1100110101",
   "111100" when "1100110110",
   "111101" when "1100110111",
   "111101" when "1100111000",
   "111101" when "1100111001",
   "111110" when "1100111010",
   "111110" when "1100111011",
   "111111" when "1100111100",
   "111111" when "1100111101",
   "111111" when "1100111110",
   "111111" when "1100111111",
   "110100" when "1101000000",
   "110100" when "1101000001",
   "110101" when "1101000010",
   "110101" when "1101000011",
   "110110" when "1101000100",
   "110110" when "1101000101",
   "110110" when "1101000110",
   "110111" when "1101000111",
   "110111" when "1101001000",
   "111000" when "1101001001",
   "111000" when "1101001010",
   "111000" when "1101001011",
   "111001" when "1101001100",
   "111001" when "1101001101",
   "111001" when "1101001110",
   "111010" when "1101001111",
   "111010" when "1101010000",
   "111011" when "1101010001",
   "111011" when "1101010010",
   "111011" when "1101010011",
   "111100" when "1101010100",
   "111100" when "1101010101",
   "111100" when "1101010110",
   "111101" when "1101010111",
   "111101" when "1101011000",
   "111110" when "1101011001",
   "111110" when "1101011010",
   "111110" when "1101011011",
   "111111" when "1101011100",
   "111111" when "1101011101",
   "111111" when "1101011110",
   "111111" when "1101011111",
   "110100" when "1101100000",
   "110101" when "1101100001",
   "110101" when "1101100010",
   "110110" when "1101100011",
   "110110" when "1101100100",
   "110110" when "1101100101",
   "110111" when "1101100110",
   "110111" when "1101100111",
   "110111" when "1101101000",
   "111000" when "1101101001",
   "111000" when "1101101010",
   "111000" when "1101101011",
   "111001" when "1101101100",
   "111001" when "1101101101",
   "111010" when "1101101110",
   "111010" when "1101101111",
   "111010" when "1101110000",
   "111011" when "1101110001",
   "111011" when "1101110010",
   "111011" when "1101110011",
   "111100" when "1101110100",
   "111100" when "1101110101",
   "111101" when "1101110110",
   "111101" when "1101110111",
   "111101" when "1101111000",
   "111110" when "1101111001",
   "111110" when "1101111010",
   "111110" when "1101111011",
   "111111" when "1101111100",
   "111111" when "1101111101",
   "111111" when "1101111110",
   "111111" when "1101111111",
   "110101" when "1110000000",
   "110101" when "1110000001",
   "110110" when "1110000010",
   "110110" when "1110000011",
   "110110" when "1110000100",
   "110111" when "1110000101",
   "110111" when "1110000110",
   "110111" when "1110000111",
   "111000" when "1110001000",
   "111000" when "1110001001",
   "111000" when "1110001010",
   "111001" when "1110001011",
   "111001" when "1110001100",
   "111001" when "1110001101",
   "111010" when "1110001110",
   "111010" when "1110001111",
   "111010" when "1110010000",
   "111011" when "1110010001",
   "111011" when "1110010010",
   "111100" when "1110010011",
   "111100" when "1110010100",
   "111100" when "1110010101",
   "111101" when "1110010110",
   "111101" when "1110010111",
   "111101" when "1110011000",
   "111110" when "1110011001",
   "111110" when "1110011010",
   "111110" when "1110011011",
   "111111" when "1110011100",
   "111111" when "1110011101",
   "111111" when "1110011110",
   "111111" when "1110011111",
   "110101" when "1110100000",
   "110110" when "1110100001",
   "110110" when "1110100010",
   "110110" when "1110100011",
   "110111" when "1110100100",
   "110111" when "1110100101",
   "110111" when "1110100110",
   "111000" when "1110100111",
   "111000" when "1110101000",
   "111000" when "1110101001",
   "111001" when "1110101010",
   "111001" when "1110101011",
   "111001" when "1110101100",
   "111010" when "1110101101",
   "111010" when "1110101110",
   "111010" when "1110101111",
   "111011" when "1110110000",
   "111011" when "1110110001",
   "111011" when "1110110010",
   "111100" when "1110110011",
   "111100" when "1110110100",
   "111100" when "1110110101",
   "111101" when "1110110110",
   "111101" when "1110110111",
   "111101" when "1110111000",
   "111110" when "1110111001",
   "111110" when "1110111010",
   "111110" when "1110111011",
   "111111" when "1110111100",
   "111111" when "1110111101",
   "111111" when "1110111110",
   "111111" when "1110111111",
   "110101" when "1111000000",
   "110110" when "1111000001",
   "110110" when "1111000010",
   "110110" when "1111000011",
   "110111" when "1111000100",
   "110111" when "1111000101",
   "110111" when "1111000110",
   "111000" when "1111000111",
   "111000" when "1111001000",
   "111000" when "1111001001",
   "111001" when "1111001010",
   "111001" when "1111001011",
   "111001" when "1111001100",
   "111010" when "1111001101",
   "111010" when "1111001110",
   "111010" when "1111001111",
   "111011" when "1111010000",
   "111011" when "1111010001",
   "111011" when "1111010010",
   "111100" when "1111010011",
   "111100" when "1111010100",
   "111100" when "1111010101",
   "111101" when "1111010110",
   "111101" when "1111010111",
   "111101" when "1111011000",
   "111110" when "1111011001",
   "111110" when "1111011010",
   "111110" when "1111011011",
   "111111" when "1111011100",
   "111111" when "1111011101",
   "111111" when "1111011110",
   "111111" when "1111011111",
   "110110" when "1111100000",
   "110110" when "1111100001",
   "110110" when "1111100010",
   "110111" when "1111100011",
   "110111" when "1111100100",
   "110111" when "1111100101",
   "111000" when "1111100110",
   "111000" when "1111100111",
   "111000" when "1111101000",
   "111001" when "1111101001",
   "111001" when "1111101010",
   "111001" when "1111101011",
   "111010" when "1111101100",
   "111010" when "1111101101",
   "111010" when "1111101110",
   "111011" when "1111101111",
   "111011" when "1111110000",
   "111011" when "1111110001",
   "111100" when "1111110010",
   "111100" when "1111110011",
   "111100" when "1111110100",
   "111101" when "1111110101",
   "111101" when "1111110110",
   "111101" when "1111110111",
   "111110" when "1111111000",
   "111110" when "1111111001",
   "111110" when "1111111010",
   "111111" when "1111111011",
   "111111" when "1111111100",
   "111111" when "1111111101",
   "111111" when "1111111110",
   "111111" when "1111111111",
   "------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                                 atan_uid36
--         (BipartiteTable_f_atan_x_pi_in_M16_out_M2_M15_F400_uid27)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Matei Istoan (2014)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity atan_uid36 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(15 downto 0);
          Y : out  std_logic_vector(13 downto 0)   );
end entity;

architecture arch of atan_uid36 is
   component GenericTable_10_16_F400_uid29 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(15 downto 0)   );
   end component;

   component GenericTable_10_6_F400_uid33 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(9 downto 0);
             Y : out  std_logic_vector(5 downto 0)   );
   end component;

signal X0 :  std_logic_vector(4 downto 0);
signal X1 :  std_logic_vector(4 downto 0);
signal X2 :  std_logic_vector(5 downto 0);
signal X2_msb :  std_logic;
signal X2_short :  std_logic_vector(4 downto 0);
signal X2_short_inv :  std_logic_vector(4 downto 0);
signal tableTIVaddr :  std_logic_vector(9 downto 0);
signal tableTOaddr :  std_logic_vector(9 downto 0);
signal tableTIVout :  std_logic_vector(15 downto 0);
signal tableTOout :  std_logic_vector(5 downto 0);
signal tableTOout_inv :  std_logic_vector(5 downto 0);
signal tableTIV_fxp :  signed(-2+17 downto 0);
signal tableTO_fxp :  signed(-12+17 downto 0);
signal tableTO_fxp_sgnExt :  signed(-2+17 downto 0);
signal Y_int :  signed(-2+17 downto 0);
signal Y_int_short :  signed(-2+16 downto 0);
signal Y_rnd :  signed(-2+16 downto 0);
attribute rom_extract: string;
attribute rom_style: string;
attribute rom_extract of GenericTable_10_16_F400_uid29: component is "yes";
attribute rom_extract of GenericTable_10_6_F400_uid33: component is "yes";
attribute rom_style of GenericTable_10_16_F400_uid29: component is "block";
attribute rom_style of GenericTable_10_6_F400_uid33: component is "block";
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   X0 <= X(15 downto 11);
   X1 <= X(10 downto 6);
   X2 <= X(5 downto 0);

   X2_msb <= X2(5);
   X2_short <= X2(4 downto 0);
   X2_short_inv <= X2_short xor (4 downto 0 => X2_msb);

   tableTIVaddr <= X0 & X1;
   tableTOaddr <= X0 & X2_short_inv;

   TIVtable: GenericTable_10_16_F400_uid29  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => tableTIVaddr,
                 Y => tableTIVout);

   TOtable: GenericTable_10_6_F400_uid33  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => tableTOaddr,
                 Y => tableTOout);

   tableTOout_inv <= tableTOout xor (5 downto 0 => X2_msb);

   tableTIV_fxp <= signed(tableTIVout);
   tableTO_fxp <= signed(tableTOout_inv);
   tableTO_fxp_sgnExt <= (9 downto 0 => tableTO_fxp(5)) & tableTO_fxp(5 downto 0); -- fix resize from (-12, -17) to (-2, -17)

   Y_int <= tableTIV_fxp + tableTO_fxp_sgnExt;
   Y_int_short <= Y_int(15 downto 1); -- fix resize from (-2, -17) to (-2, -16)
   Y_rnd <= Y_int_short + ("00000000000000" & '1');
   Y <= std_logic_vector(Y_rnd(14 downto 1));
end architecture;

--------------------------------------------------------------------------------
--                  FixAtan2ByRecipMultAtan_16_16_F400_uid2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Matei Istoan, Florent de Dinechin (2012-...)
--------------------------------------------------------------------------------
-- Pipeline depth: 5 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixAtan2ByRecipMultAtan_16_16_F400_uid2 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(15 downto 0);
          Y : in  std_logic_vector(15 downto 0);
          A : out  std_logic_vector(15 downto 0)   );
end entity;

architecture arch of FixAtan2ByRecipMultAtan_16_16_F400_uid2 is
   component LZOC_14_F400_uid4 is
      port ( clk, rst : in std_logic;
             I : in  std_logic_vector(13 downto 0);
             OZB : in  std_logic;
             O : out  std_logic_vector(3 downto 0)   );
   end component;

   component LeftShifter_15_by_max_14_F400_uid8 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(14 downto 0);
             S : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(28 downto 0)   );
   end component;

   component reciprocal_uid23 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(13 downto 0);
             Y : out  std_logic_vector(17 downto 0)   );
   end component;

   component atan_uid36 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(15 downto 0);
             Y : out  std_logic_vector(13 downto 0)   );
   end component;

signal sgnX :  std_logic;
signal sgnY :  std_logic;
signal Xsat :  std_logic_vector(15 downto 0);
signal Ysat :  std_logic_vector(15 downto 0);
signal pX :  std_logic_vector(15 downto 0);
signal pY :  std_logic_vector(15 downto 0);
signal mX :  std_logic_vector(15 downto 0);
signal mY :  std_logic_vector(15 downto 0);
signal XmY :  std_logic_vector(16 downto 0);
signal XpY :  std_logic_vector(16 downto 0);
signal XltY :  std_logic;
signal mYltX :  std_logic;
signal quadrant, quadrant_d1, quadrant_d2, quadrant_d3, quadrant_d4, quadrant_d5 :  std_logic_vector(1 downto 0);
signal XR, XR_d1, XR_d2, XR_d3 :  std_logic_vector(14 downto 0);
signal YR, YR_d1, YR_d2, YR_d3 :  std_logic_vector(14 downto 0);
signal finalAdd, finalAdd_d1, finalAdd_d2, finalAdd_d3, finalAdd_d4, finalAdd_d5 :  std_logic;
signal XorY :  std_logic_vector(13 downto 0);
signal S :  std_logic_vector(3 downto 0);
signal XRSfull :  std_logic_vector(28 downto 0);
signal XRS, XRS_d1 :  std_logic_vector(14 downto 0);
signal YRSfull :  std_logic_vector(28 downto 0);
signal YRS, YRS_d1 :  std_logic_vector(14 downto 0);
signal XRm1 :  std_logic_vector(13 downto 0);
signal R0 :  std_logic_vector(17 downto 0);
signal R, R_d1 :  unsigned(0+16 downto 0);
signal YRU, YRU_d1 :  unsigned(-1+15 downto 0);
signal P :  unsigned(0+31 downto 0);
signal PtruncU :  unsigned(-1+16 downto 0);
signal P_slv :  std_logic_vector(15 downto 0);
signal atanTableOut :  std_logic_vector(13 downto 0);
signal finalZ :  std_logic_vector(15 downto 0);
signal qangle :  std_logic_vector(15 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            quadrant_d1 <=  quadrant;
            quadrant_d2 <=  quadrant_d1;
            quadrant_d3 <=  quadrant_d2;
            quadrant_d4 <=  quadrant_d3;
            quadrant_d5 <=  quadrant_d4;
            XR_d1 <=  XR;
            XR_d2 <=  XR_d1;
            XR_d3 <=  XR_d2;
            YR_d1 <=  YR;
            YR_d2 <=  YR_d1;
            YR_d3 <=  YR_d2;
            finalAdd_d1 <=  finalAdd;
            finalAdd_d2 <=  finalAdd_d1;
            finalAdd_d3 <=  finalAdd_d2;
            finalAdd_d4 <=  finalAdd_d3;
            finalAdd_d5 <=  finalAdd_d4;
            XRS_d1 <=  XRS;
            YRS_d1 <=  YRS;
            R_d1 <=  R;
            YRU_d1 <=  YRU;
         end if;
      end process;
   sgnX <= X(15);
   sgnY <= Y(15);
   -- First saturate x and y in case they touch -1
   Xsat <= "1000000000000001" when X="1000000000000000" else X ;
   Ysat <= "1000000000000001" when Y="1000000000000000" else Y ;
   pX <= Xsat;
   pY <= Ysat;
   mX <= ("0000000000000000" - Xsat);
   mY <= ("0000000000000000" - Ysat);
   XmY <= (sgnX & Xsat)-(sgnY & Ysat);
   XpY <= (sgnX & Xsat)+(sgnY & Ysat);
   XltY <= XmY(16);
   mYltX <= not XpY(16);
   -- quadrant will also be the angle to add at the end
   quadrant <= 
      "00"  when (not sgnX and not XltY and     mYltX)='1' else
      "01"  when (not sgnY and     XltY and     mYltX)='1' else
      "10"  when (    sgnX and     XltY and not mYltX)='1' else
      "11";
   XR <= 
      pX(14 downto 0) when quadrant="00"   else 
      pY(14 downto 0) when quadrant="01"   else 
      mX(14 downto 0) when quadrant="10"   else 
      mY(14 downto 0);
   YR <= 
      pY(14 downto 0) when quadrant="00" and sgnY='0'  else 
      mY(14 downto 0) when quadrant="00" and sgnY='1'  else 
      pX(14 downto 0) when quadrant="01" and sgnX='0'  else 
      mX(14 downto 0) when quadrant="01" and sgnX='1'  else 
      pY(14 downto 0) when quadrant="10" and sgnY='0'  else 
      mY(14 downto 0) when quadrant="10" and sgnY='1'  else 
      pX(14 downto 0) when quadrant="11" and sgnX='0'  else 
      mX(14 downto 0) ;
   finalAdd <= 
      '1' when (quadrant="00" and sgnY='0') or(quadrant="01" and sgnX='1') or (quadrant="10" and sgnY='1') or (quadrant="11" and sgnX='0')
       else '0';  -- this information is sent to the end of the pipeline, better compute it here as one bit
   ----------------Synchro barrier, entering cycle 1----------------
   XorY <= XR_d1(14 downto 1) or YR_d1(14 downto 1);
   lzc: LZOC_14_F400_uid4  -- pipelineDepth=2 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 I => XorY,
                 O => S,
                 OZB => '0');
   ----------------Synchro barrier, entering cycle 3----------------
   Xshift: LeftShifter_15_by_max_14_F400_uid8  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => XRSfull,
                 S => S,
                 X => XR_d3);
   XRS <=  XRSfull (14 downto 0);
   Yshift: LeftShifter_15_by_max_14_F400_uid8  -- pipelineDepth=1 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 R => YRSfull,
                 S => S,
                 X => YR_d3);
   YRS <=  YRSfull (14 downto 0);
   ----------------Synchro barrier, entering cycle 4----------------
   XRm1 <= XRS_d1(13 downto 0); -- removing the MSB which is constantly 1
   recipTable: reciprocal_uid23  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => XRm1,
                 Y => R0);
   R <= unsigned(R0(16 downto 0)); -- removing the sign  bit
   YRU <= unsigned(YRS_d1);
   ----------------Synchro barrier, entering cycle 5----------------
   P <= R_d1*YRU_d1;
   PtruncU <= P(30 downto 15); -- fix resize from (0, -31) to (-1, -16)
   P_slv <=  std_logic_vector(PtruncU);
   atanTable: atan_uid36  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => P_slv,
                 Y => atanTableOut);
   finalZ <= "00" & atanTableOut;
   qangle <= (quadrant_d5 & "00000000000000");
   A <=            qangle + finalZ  when finalAdd_d5='1'
      else qangle - finalZ;
end architecture;

