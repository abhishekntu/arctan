--------------------------------------------------------------------------------
--                             LZOC_12_F400_uid4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- Pipeline depth: 2 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOC_12_F400_uid4 is
   port ( clk, rst : in std_logic;
          I : in  std_logic_vector(11 downto 0);
          OZB : in  std_logic;
          O : out  std_logic_vector(3 downto 0)   );
end entity;

architecture arch of LZOC_12_F400_uid4 is
signal sozb, sozb_d1, sozb_d2 :  std_logic;
signal level4, level4_d1 :  std_logic_vector(15 downto 0);
signal digit4, digit4_d1 :  std_logic;
signal level3 :  std_logic_vector(7 downto 0);
signal digit3, digit3_d1 :  std_logic;
signal level2, level2_d1 :  std_logic_vector(3 downto 0);
signal digit2 :  std_logic;
signal level1 :  std_logic_vector(1 downto 0);
signal digit1 :  std_logic;
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            sozb_d1 <=  sozb;
            sozb_d2 <=  sozb_d1;
            level4_d1 <=  level4;
            digit4_d1 <=  digit4;
            digit3_d1 <=  digit3;
            level2_d1 <=  level2;
         end if;
      end process;
   sozb <= OZB;
   level4<= I& (3 downto 0 => not(sozb));
   ----------------Synchro barrier, entering cycle 1----------------
   digit4<= '1' when level4_d1(15 downto 8) = (15 downto 8 => sozb_d1) else '0';
   level3<= level4_d1(7 downto 0) when digit4='1' else level4_d1(15 downto 8);
   digit3<= '1' when level3(7 downto 4) = (7 downto 4 => sozb_d1) else '0';
   level2<= level3(3 downto 0) when digit3='1' else level3(7 downto 4);
   ----------------Synchro barrier, entering cycle 2----------------
   digit2<= '1' when level2_d1(3 downto 2) = (3 downto 2 => sozb_d2) else '0';
   level1<= level2_d1(1 downto 0) when digit2='1' else level2_d1(3 downto 2);
   digit1<= '1' when level1(1 downto 1) = (1 downto 1 => sozb_d2) else '0';
   O <= digit4_d1 & digit3_d1 & digit2 & digit1;
end architecture;

--------------------------------------------------------------------------------
--                     LeftShifter_13_by_max_12_F400_uid8
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- Pipeline depth: 1 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter_13_by_max_12_F400_uid8 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(12 downto 0);
          S : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(24 downto 0)   );
end entity;

architecture arch of LeftShifter_13_by_max_12_F400_uid8 is
signal level0 :  std_logic_vector(12 downto 0);
signal ps, ps_d1 :  std_logic_vector(3 downto 0);
signal level1 :  std_logic_vector(13 downto 0);
signal level2 :  std_logic_vector(15 downto 0);
signal level3, level3_d1 :  std_logic_vector(19 downto 0);
signal level4 :  std_logic_vector(27 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            ps_d1 <=  ps;
            level3_d1 <=  level3;
         end if;
      end process;
   level0<= X;
   ps<= S;
   level1<= level0 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => '0') & level0;
   level2<= level1 & (1 downto 0 => '0') when ps(1)= '1' else     (1 downto 0 => '0') & level1;
   level3<= level2 & (3 downto 0 => '0') when ps(2)= '1' else     (3 downto 0 => '0') & level2;
   ----------------Synchro barrier, entering cycle 1----------------
   level4<= level3_d1 & (7 downto 0 => '0') when ps_d1(3)= '1' else     (7 downto 0 => '0') & level3_d1;
   R <= level4(24 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                        GenericTable_8_18_F400_uid16
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity GenericTable_8_18_F400_uid16 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          Y : out  std_logic_vector(17 downto 0)   );
end entity;

architecture arch of GenericTable_8_18_F400_uid16 is
signal TableOut :  std_logic_vector(17 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
  with X select TableOut <= 
   "011111111100001101" when "00000000",
   "011111110100010001" when "00000001",
   "011111101100011001" when "00000010",
   "011111100100100100" when "00000011",
   "011111011100110100" when "00000100",
   "011111010101000111" when "00000101",
   "011111001101011110" when "00000110",
   "011111000101111001" when "00000111",
   "011110111110010111" when "00001000",
   "011110110110111001" when "00001001",
   "011110101111011111" when "00001010",
   "011110101000001000" when "00001011",
   "011110100000110101" when "00001100",
   "011110011001100101" when "00001101",
   "011110010010011001" when "00001110",
   "011110001011010000" when "00001111",
   "011110000100001010" when "00010000",
   "011101111101001000" when "00010001",
   "011101110110001001" when "00010010",
   "011101101111001101" when "00010011",
   "011101101000010100" when "00010100",
   "011101100001011111" when "00010101",
   "011101011010101101" when "00010110",
   "011101010011111101" when "00010111",
   "011101001101010001" when "00011000",
   "011101000110101000" when "00011001",
   "011101000000000010" when "00011010",
   "011100111001011111" when "00011011",
   "011100110010111111" when "00011100",
   "011100101100100010" when "00011101",
   "011100100110000111" when "00011110",
   "011100011111110000" when "00011111",
   "011100011001011011" when "00100000",
   "011100010011001010" when "00100001",
   "011100001100111011" when "00100010",
   "011100000110101110" when "00100011",
   "011100000000100101" when "00100100",
   "011011111010011110" when "00100101",
   "011011110100011001" when "00100110",
   "011011101110011000" when "00100111",
   "011011101000011001" when "00101000",
   "011011100010011100" when "00101001",
   "011011011100100010" when "00101010",
   "011011010110101011" when "00101011",
   "011011010000110110" when "00101100",
   "011011001011000011" when "00101101",
   "011011000101010011" when "00101110",
   "011010111111100110" when "00101111",
   "011010111001111011" when "00110000",
   "011010110100010010" when "00110001",
   "011010101110101100" when "00110010",
   "011010101001000111" when "00110011",
   "011010100011100110" when "00110100",
   "011010011110000110" when "00110101",
   "011010011000101001" when "00110110",
   "011010010011001110" when "00110111",
   "011010001101110101" when "00111000",
   "011010001000011111" when "00111001",
   "011010000011001010" when "00111010",
   "011001111101111000" when "00111011",
   "011001111000101000" when "00111100",
   "011001110011011010" when "00111101",
   "011001101110001110" when "00111110",
   "011001101001000100" when "00111111",
   "011001100011111100" when "01000000",
   "011001011110110111" when "01000001",
   "011001011001110011" when "01000010",
   "011001010100110001" when "01000011",
   "011001001111110010" when "01000100",
   "011001001010110100" when "01000101",
   "011001000101111000" when "01000110",
   "011001000000111110" when "01000111",
   "011000111100000110" when "01001000",
   "011000110111010000" when "01001001",
   "011000110010011100" when "01001010",
   "011000101101101010" when "01001011",
   "011000101000111001" when "01001100",
   "011000100100001011" when "01001101",
   "011000011111011110" when "01001110",
   "011000011010110011" when "01001111",
   "011000010110001001" when "01010000",
   "011000010001100010" when "01010001",
   "011000001100111100" when "01010010",
   "011000001000011000" when "01010011",
   "011000000011110110" when "01010100",
   "010111111111010101" when "01010101",
   "010111111010110110" when "01010110",
   "010111110110011001" when "01010111",
   "010111110001111101" when "01011000",
   "010111101101100011" when "01011001",
   "010111101001001011" when "01011010",
   "010111100100110100" when "01011011",
   "010111100000011111" when "01011100",
   "010111011100001100" when "01011101",
   "010111010111111010" when "01011110",
   "010111010011101001" when "01011111",
   "010111001111011010" when "01100000",
   "010111001011001101" when "01100001",
   "010111000111000001" when "01100010",
   "010111000010110111" when "01100011",
   "010110111110101110" when "01100100",
   "010110111010100111" when "01100101",
   "010110110110100001" when "01100110",
   "010110110010011101" when "01100111",
   "010110101110011010" when "01101000",
   "010110101010011000" when "01101001",
   "010110100110011000" when "01101010",
   "010110100010011001" when "01101011",
   "010110011110011100" when "01101100",
   "010110011010100000" when "01101101",
   "010110010110100110" when "01101110",
   "010110010010101100" when "01101111",
   "010110001110110101" when "01110000",
   "010110001010111110" when "01110001",
   "010110000111001001" when "01110010",
   "010110000011010101" when "01110011",
   "010101111111100011" when "01110100",
   "010101111011110010" when "01110101",
   "010101111000000010" when "01110110",
   "010101110100010011" when "01110111",
   "010101110000100110" when "01111000",
   "010101101100111001" when "01111001",
   "010101101001001111" when "01111010",
   "010101100101100101" when "01111011",
   "010101100001111100" when "01111100",
   "010101011110010101" when "01111101",
   "010101011010101111" when "01111110",
   "010101010111001011" when "01111111",
   "010101010011100111" when "10000000",
   "010101010000000101" when "10000001",
   "010101001100100011" when "10000010",
   "010101001001000011" when "10000011",
   "010101000101100100" when "10000100",
   "010101000010000111" when "10000101",
   "010100111110101010" when "10000110",
   "010100111011001110" when "10000111",
   "010100110111110100" when "10001000",
   "010100110100011011" when "10001001",
   "010100110001000010" when "10001010",
   "010100101101101011" when "10001011",
   "010100101010010101" when "10001100",
   "010100100111000000" when "10001101",
   "010100100011101101" when "10001110",
   "010100100000011010" when "10001111",
   "010100011101001000" when "10010000",
   "010100011001110111" when "10010001",
   "010100010110101000" when "10010010",
   "010100010011011001" when "10010011",
   "010100010000001011" when "10010100",
   "010100001100111111" when "10010101",
   "010100001001110011" when "10010110",
   "010100000110101001" when "10010111",
   "010100000011011111" when "10011000",
   "010100000000010110" when "10011001",
   "010011111101001111" when "10011010",
   "010011111010001000" when "10011011",
   "010011110111000010" when "10011100",
   "010011110011111110" when "10011101",
   "010011110000111010" when "10011110",
   "010011101101110111" when "10011111",
   "010011101010110101" when "10100000",
   "010011100111110100" when "10100001",
   "010011100100110100" when "10100010",
   "010011100001110101" when "10100011",
   "010011011110110111" when "10100100",
   "010011011011111001" when "10100101",
   "010011011000111101" when "10100110",
   "010011010110000001" when "10100111",
   "010011010011000111" when "10101000",
   "010011010000001101" when "10101001",
   "010011001101010100" when "10101010",
   "010011001010011100" when "10101011",
   "010011000111100101" when "10101100",
   "010011000100101110" when "10101101",
   "010011000001111001" when "10101110",
   "010010111111000100" when "10101111",
   "010010111100010000" when "10110000",
   "010010111001011101" when "10110001",
   "010010110110101011" when "10110010",
   "010010110011111010" when "10110011",
   "010010110001001001" when "10110100",
   "010010101110011001" when "10110101",
   "010010101011101010" when "10110110",
   "010010101000111100" when "10110111",
   "010010100110001111" when "10111000",
   "010010100011100010" when "10111001",
   "010010100000110111" when "10111010",
   "010010011110001100" when "10111011",
   "010010011011100001" when "10111100",
   "010010011000111000" when "10111101",
   "010010010110001111" when "10111110",
   "010010010011100111" when "10111111",
   "010010010001000000" when "11000000",
   "010010001110011010" when "11000001",
   "010010001011110100" when "11000010",
   "010010001001001111" when "11000011",
   "010010000110101011" when "11000100",
   "010010000100000111" when "11000101",
   "010010000001100100" when "11000110",
   "010001111111000010" when "11000111",
   "010001111100100001" when "11001000",
   "010001111010000000" when "11001001",
   "010001110111100000" when "11001010",
   "010001110101000001" when "11001011",
   "010001110010100010" when "11001100",
   "010001110000000100" when "11001101",
   "010001101101100111" when "11001110",
   "010001101011001011" when "11001111",
   "010001101000101111" when "11010000",
   "010001100110010011" when "11010001",
   "010001100011111001" when "11010010",
   "010001100001011111" when "11010011",
   "010001011111000110" when "11010100",
   "010001011100101101" when "11010101",
   "010001011010010101" when "11010110",
   "010001010111111110" when "11010111",
   "010001010101100111" when "11011000",
   "010001010011010001" when "11011001",
   "010001010000111100" when "11011010",
   "010001001110100111" when "11011011",
   "010001001100010011" when "11011100",
   "010001001010000000" when "11011101",
   "010001000111101101" when "11011110",
   "010001000101011011" when "11011111",
   "010001000011001001" when "11100000",
   "010001000000111000" when "11100001",
   "010000111110100111" when "11100010",
   "010000111100011000" when "11100011",
   "010000111010001000" when "11100100",
   "010000110111111010" when "11100101",
   "010000110101101100" when "11100110",
   "010000110011011110" when "11100111",
   "010000110001010001" when "11101000",
   "010000101111000101" when "11101001",
   "010000101100111001" when "11101010",
   "010000101010101110" when "11101011",
   "010000101000100011" when "11101100",
   "010000100110011001" when "11101101",
   "010000100100010000" when "11101110",
   "010000100010000111" when "11101111",
   "010000011111111110" when "11110000",
   "010000011101110110" when "11110001",
   "010000011011101111" when "11110010",
   "010000011001101000" when "11110011",
   "010000010111100010" when "11110100",
   "010000010101011100" when "11110101",
   "010000010011010111" when "11110110",
   "010000010001010011" when "11110111",
   "010000001111001110" when "11111000",
   "010000001101001011" when "11111001",
   "010000001011001000" when "11111010",
   "010000001001000101" when "11111011",
   "010000000111000011" when "11111100",
   "010000000101000010" when "11111101",
   "010000000011000001" when "11111110",
   "010000000001000000" when "11111111",
   "------------------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                        GenericTable_7_10_F400_uid20
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity GenericTable_7_10_F400_uid20 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(6 downto 0);
          Y : out  std_logic_vector(9 downto 0)   );
end entity;

architecture arch of GenericTable_7_10_F400_uid20 is
signal TableOut :  std_logic_vector(9 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
  with X select TableOut <= 
   "0011100010" when "0000000",
   "0011000100" when "0000001",
   "0010100110" when "0000010",
   "0010000111" when "0000011",
   "0001101001" when "0000100",
   "0001001011" when "0000101",
   "0000101101" when "0000110",
   "0000001111" when "0000111",
   "0011001001" when "0001000",
   "0010101110" when "0001001",
   "0010010011" when "0001010",
   "0001111000" when "0001011",
   "0001011110" when "0001100",
   "0001000011" when "0001101",
   "0000101000" when "0001110",
   "0000001101" when "0001111",
   "0010110100" when "0010000",
   "0010011100" when "0010001",
   "0010000100" when "0010010",
   "0001101100" when "0010011",
   "0001010100" when "0010100",
   "0000111100" when "0010101",
   "0000100100" when "0010110",
   "0000001100" when "0010111",
   "0010100010" when "0011000",
   "0010001100" when "0011001",
   "0001110111" when "0011010",
   "0001100001" when "0011011",
   "0001001011" when "0011100",
   "0000110110" when "0011101",
   "0000100000" when "0011110",
   "0000001011" when "0011111",
   "0010010010" when "0100000",
   "0001111111" when "0100001",
   "0001101011" when "0100010",
   "0001011000" when "0100011",
   "0001000100" when "0100100",
   "0000110001" when "0100101",
   "0000011101" when "0100110",
   "0000001010" when "0100111",
   "0010000101" when "0101000",
   "0001110011" when "0101001",
   "0001100001" when "0101010",
   "0001010000" when "0101011",
   "0000111110" when "0101100",
   "0000101100" when "0101101",
   "0000011011" when "0101110",
   "0000001001" when "0101111",
   "0001111001" when "0110000",
   "0001101001" when "0110001",
   "0001011001" when "0110010",
   "0001001001" when "0110011",
   "0000111001" when "0110100",
   "0000101000" when "0110101",
   "0000011000" when "0110110",
   "0000001000" when "0110111",
   "0001101111" when "0111000",
   "0001100000" when "0111001",
   "0001010010" when "0111010",
   "0001000011" when "0111011",
   "0000110100" when "0111100",
   "0000100101" when "0111101",
   "0000010110" when "0111110",
   "0000000111" when "0111111",
   "0001100110" when "1000000",
   "0001011001" when "1000001",
   "0001001011" when "1000010",
   "0000111101" when "1000011",
   "0000110000" when "1000100",
   "0000100010" when "1000101",
   "0000010100" when "1000110",
   "0000000111" when "1000111",
   "0001011111" when "1001000",
   "0001010010" when "1001001",
   "0001000101" when "1001010",
   "0000111001" when "1001011",
   "0000101100" when "1001100",
   "0000100000" when "1001101",
   "0000010011" when "1001110",
   "0000000110" when "1001111",
   "0001011000" when "1010000",
   "0001001100" when "1010001",
   "0001000000" when "1010010",
   "0000110101" when "1010011",
   "0000101001" when "1010100",
   "0000011101" when "1010101",
   "0000010010" when "1010110",
   "0000000110" when "1010111",
   "0001010001" when "1011000",
   "0001000110" when "1011001",
   "0000111100" when "1011010",
   "0000110001" when "1011011",
   "0000100110" when "1011100",
   "0000011011" when "1011101",
   "0000010000" when "1011110",
   "0000000101" when "1011111",
   "0001001100" when "1100000",
   "0001000010" when "1100001",
   "0000110111" when "1100010",
   "0000101101" when "1100011",
   "0000100011" when "1100100",
   "0000011001" when "1100101",
   "0000001111" when "1100110",
   "0000000101" when "1100111",
   "0001000111" when "1101000",
   "0000111101" when "1101001",
   "0000110100" when "1101010",
   "0000101010" when "1101011",
   "0000100001" when "1101100",
   "0000011000" when "1101101",
   "0000001110" when "1101110",
   "0000000101" when "1101111",
   "0001000010" when "1110000",
   "0000111001" when "1110001",
   "0000110000" when "1110010",
   "0000101000" when "1110011",
   "0000011111" when "1110100",
   "0000010110" when "1110101",
   "0000001101" when "1110110",
   "0000000100" when "1110111",
   "0000111110" when "1111000",
   "0000110110" when "1111001",
   "0000101101" when "1111010",
   "0000100101" when "1111011",
   "0000011101" when "1111100",
   "0000010101" when "1111101",
   "0000001100" when "1111110",
   "0000000100" when "1111111",
   "----------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                              reciprocal_uid23
--        (BipartiteTable_f_2_1Px_M1bM14_in_M12_out_1_M14_F400_uid14)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Matei Istoan (2014)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity reciprocal_uid23 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(11 downto 0);
          Y : out  std_logic_vector(15 downto 0)   );
end entity;

architecture arch of reciprocal_uid23 is
   component GenericTable_8_18_F400_uid16 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             Y : out  std_logic_vector(17 downto 0)   );
   end component;

   component GenericTable_7_10_F400_uid20 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(6 downto 0);
             Y : out  std_logic_vector(9 downto 0)   );
   end component;

signal X0 :  std_logic_vector(3 downto 0);
signal X1 :  std_logic_vector(3 downto 0);
signal X2 :  std_logic_vector(3 downto 0);
signal X2_msb :  std_logic;
signal X2_short :  std_logic_vector(2 downto 0);
signal X2_short_inv :  std_logic_vector(2 downto 0);
signal tableTIVaddr :  std_logic_vector(7 downto 0);
signal tableTOaddr :  std_logic_vector(6 downto 0);
signal tableTIVout :  std_logic_vector(17 downto 0);
signal tableTOout :  std_logic_vector(9 downto 0);
signal tableTOout_inv :  std_logic_vector(9 downto 0);
signal tableTIV_fxp :  signed(1+16 downto 0);
signal tableTO_fxp :  signed(-7+16 downto 0);
signal tableTO_fxp_sgnExt :  signed(1+16 downto 0);
signal Y_int :  signed(1+16 downto 0);
signal Y_int_short :  signed(1+15 downto 0);
signal Y_rnd :  signed(1+15 downto 0);
attribute rom_extract: string;
attribute rom_style: string;
attribute rom_extract of GenericTable_7_10_F400_uid20: component is "yes";
attribute rom_extract of GenericTable_8_18_F400_uid16: component is "yes";
attribute rom_style of GenericTable_7_10_F400_uid20: component is "block";
attribute rom_style of GenericTable_8_18_F400_uid16: component is "block";
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   X0 <= X(11 downto 8);
   X1 <= X(7 downto 4);
   X2 <= X(3 downto 0);

   X2_msb <= X2(3);
   X2_short <= X2(2 downto 0);
   X2_short_inv <= X2_short xor (2 downto 0 => X2_msb);

   tableTIVaddr <= X0 & X1;
   tableTOaddr <= X0 & X2_short_inv;

   TIVtable: GenericTable_8_18_F400_uid16  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => tableTIVaddr,
                 Y => tableTIVout);

   TOtable: GenericTable_7_10_F400_uid20  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => tableTOaddr,
                 Y => tableTOout);

   tableTOout_inv <= tableTOout xor (9 downto 0 => X2_msb);

   tableTIV_fxp <= signed(tableTIVout);
   tableTO_fxp <= signed(tableTOout_inv);
   tableTO_fxp_sgnExt <= (7 downto 0 => tableTO_fxp(9)) & tableTO_fxp(9 downto 0); -- fix resize from (-7, -16) to (1, -16)

   Y_int <= tableTIV_fxp + tableTO_fxp_sgnExt;
   Y_int_short <= Y_int(17 downto 1); -- fix resize from (1, -16) to (1, -15)
   Y_rnd <= Y_int_short + ("0000000000000000" & '1');
   Y <= std_logic_vector(Y_rnd(16 downto 1));
end architecture;

--------------------------------------------------------------------------------
--                        GenericTable_8_14_F400_uid29
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity GenericTable_8_14_F400_uid29 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(7 downto 0);
          Y : out  std_logic_vector(13 downto 0)   );
end entity;

architecture arch of GenericTable_8_14_F400_uid29 is
signal TableOut :  std_logic_vector(13 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
  with X select TableOut <= 
   "00000000010100" when "00000000",
   "00000000111101" when "00000001",
   "00000001100110" when "00000010",
   "00000010001110" when "00000011",
   "00000010110111" when "00000100",
   "00000011100000" when "00000101",
   "00000100001000" when "00000110",
   "00000100110001" when "00000111",
   "00000101011010" when "00001000",
   "00000110000011" when "00001001",
   "00000110101011" when "00001010",
   "00000111010100" when "00001011",
   "00000111111101" when "00001100",
   "00001000100101" when "00001101",
   "00001001001110" when "00001110",
   "00001001110110" when "00001111",
   "00001010011111" when "00010000",
   "00001011001000" when "00010001",
   "00001011110000" when "00010010",
   "00001100011001" when "00010011",
   "00001101000001" when "00010100",
   "00001101101010" when "00010101",
   "00001110010010" when "00010110",
   "00001110111010" when "00010111",
   "00001111100011" when "00011000",
   "00010000001011" when "00011001",
   "00010000110100" when "00011010",
   "00010001011100" when "00011011",
   "00010010000100" when "00011100",
   "00010010101100" when "00011101",
   "00010011010101" when "00011110",
   "00010011111101" when "00011111",
   "00010100100101" when "00100000",
   "00010101001101" when "00100001",
   "00010101110101" when "00100010",
   "00010110011101" when "00100011",
   "00010111000101" when "00100100",
   "00010111101101" when "00100101",
   "00011000010101" when "00100110",
   "00011000111100" when "00100111",
   "00011001100100" when "00101000",
   "00011010001100" when "00101001",
   "00011010110100" when "00101010",
   "00011011011011" when "00101011",
   "00011100000011" when "00101100",
   "00011100101010" when "00101101",
   "00011101010010" when "00101110",
   "00011101111001" when "00101111",
   "00011110100001" when "00110000",
   "00011111001000" when "00110001",
   "00011111101111" when "00110010",
   "00100000010110" when "00110011",
   "00100000111101" when "00110100",
   "00100001100101" when "00110101",
   "00100010001100" when "00110110",
   "00100010110011" when "00110111",
   "00100011011001" when "00111000",
   "00100100000000" when "00111001",
   "00100100100111" when "00111010",
   "00100101001110" when "00111011",
   "00100101110100" when "00111100",
   "00100110011011" when "00111101",
   "00100111000001" when "00111110",
   "00100111101000" when "00111111",
   "00101000001110" when "01000000",
   "00101000110100" when "01000001",
   "00101001011011" when "01000010",
   "00101010000001" when "01000011",
   "00101010100111" when "01000100",
   "00101011001101" when "01000101",
   "00101011110011" when "01000110",
   "00101100011000" when "01000111",
   "00101100111110" when "01001000",
   "00101101100100" when "01001001",
   "00101110001010" when "01001010",
   "00101110101111" when "01001011",
   "00101111010100" when "01001100",
   "00101111111010" when "01001101",
   "00110000011111" when "01001110",
   "00110001000100" when "01001111",
   "00110001101001" when "01010000",
   "00110010001110" when "01010001",
   "00110010110011" when "01010010",
   "00110011011000" when "01010011",
   "00110011111101" when "01010100",
   "00110100100010" when "01010101",
   "00110101000110" when "01010110",
   "00110101101011" when "01010111",
   "00110110001111" when "01011000",
   "00110110110100" when "01011001",
   "00110111011000" when "01011010",
   "00110111111100" when "01011011",
   "00111000100000" when "01011100",
   "00111001000100" when "01011101",
   "00111001101000" when "01011110",
   "00111010001100" when "01011111",
   "00111010110000" when "01100000",
   "00111011010011" when "01100001",
   "00111011110111" when "01100010",
   "00111100011010" when "01100011",
   "00111100111110" when "01100100",
   "00111101100001" when "01100101",
   "00111110000100" when "01100110",
   "00111110100111" when "01100111",
   "00111111001010" when "01101000",
   "00111111101101" when "01101001",
   "01000000010000" when "01101010",
   "01000000110010" when "01101011",
   "01000001010101" when "01101100",
   "01000001111000" when "01101101",
   "01000010011010" when "01101110",
   "01000010111100" when "01101111",
   "01000011011110" when "01110000",
   "01000100000001" when "01110001",
   "01000100100011" when "01110010",
   "01000101000100" when "01110011",
   "01000101100110" when "01110100",
   "01000110001000" when "01110101",
   "01000110101010" when "01110110",
   "01000111001011" when "01110111",
   "01000111101100" when "01111000",
   "01001000001110" when "01111001",
   "01001000101111" when "01111010",
   "01001001010000" when "01111011",
   "01001001110001" when "01111100",
   "01001010010010" when "01111101",
   "01001010110011" when "01111110",
   "01001011010011" when "01111111",
   "01001011110100" when "10000000",
   "01001100010101" when "10000001",
   "01001100110101" when "10000010",
   "01001101010101" when "10000011",
   "01001101110101" when "10000100",
   "01001110010101" when "10000101",
   "01001110110101" when "10000110",
   "01001111010101" when "10000111",
   "01001111110101" when "10001000",
   "01010000010101" when "10001001",
   "01010000110100" when "10001010",
   "01010001010100" when "10001011",
   "01010001110011" when "10001100",
   "01010010010010" when "10001101",
   "01010010110010" when "10001110",
   "01010011010001" when "10001111",
   "01010011110000" when "10010000",
   "01010100001110" when "10010001",
   "01010100101101" when "10010010",
   "01010101001100" when "10010011",
   "01010101101010" when "10010100",
   "01010110001001" when "10010101",
   "01010110100111" when "10010110",
   "01010111000101" when "10010111",
   "01010111100100" when "10011000",
   "01011000000010" when "10011001",
   "01011000011111" when "10011010",
   "01011000111101" when "10011011",
   "01011001011011" when "10011100",
   "01011001111001" when "10011101",
   "01011010010110" when "10011110",
   "01011010110011" when "10011111",
   "01011011010001" when "10100000",
   "01011011101110" when "10100001",
   "01011100001011" when "10100010",
   "01011100101000" when "10100011",
   "01011101000101" when "10100100",
   "01011101100010" when "10100101",
   "01011101111110" when "10100110",
   "01011110011011" when "10100111",
   "01011110110111" when "10101000",
   "01011111010100" when "10101001",
   "01011111110000" when "10101010",
   "01100000001100" when "10101011",
   "01100000101000" when "10101100",
   "01100001000100" when "10101101",
   "01100001100000" when "10101110",
   "01100001111100" when "10101111",
   "01100010011000" when "10110000",
   "01100010110011" when "10110001",
   "01100011001111" when "10110010",
   "01100011101010" when "10110011",
   "01100100000101" when "10110100",
   "01100100100001" when "10110101",
   "01100100111100" when "10110110",
   "01100101010111" when "10110111",
   "01100101110001" when "10111000",
   "01100110001100" when "10111001",
   "01100110100111" when "10111010",
   "01100111000001" when "10111011",
   "01100111011100" when "10111100",
   "01100111110110" when "10111101",
   "01101000010001" when "10111110",
   "01101000101011" when "10111111",
   "01101001000101" when "11000000",
   "01101001011111" when "11000001",
   "01101001111001" when "11000010",
   "01101010010010" when "11000011",
   "01101010101100" when "11000100",
   "01101011000110" when "11000101",
   "01101011011111" when "11000110",
   "01101011111001" when "11000111",
   "01101100010010" when "11001000",
   "01101100101011" when "11001001",
   "01101101000100" when "11001010",
   "01101101011101" when "11001011",
   "01101101110110" when "11001100",
   "01101110001111" when "11001101",
   "01101110101000" when "11001110",
   "01101111000000" when "11001111",
   "01101111011001" when "11010000",
   "01101111110001" when "11010001",
   "01110000001010" when "11010010",
   "01110000100010" when "11010011",
   "01110000111010" when "11010100",
   "01110001010010" when "11010101",
   "01110001101010" when "11010110",
   "01110010000010" when "11010111",
   "01110010011010" when "11011000",
   "01110010110010" when "11011001",
   "01110011001001" when "11011010",
   "01110011100001" when "11011011",
   "01110011111000" when "11011100",
   "01110100010000" when "11011101",
   "01110100100111" when "11011110",
   "01110100111110" when "11011111",
   "01110101010101" when "11100000",
   "01110101101100" when "11100001",
   "01110110000011" when "11100010",
   "01110110011010" when "11100011",
   "01110110110000" when "11100100",
   "01110111000111" when "11100101",
   "01110111011110" when "11100110",
   "01110111110100" when "11100111",
   "01111000001010" when "11101000",
   "01111000100001" when "11101001",
   "01111000110111" when "11101010",
   "01111001001101" when "11101011",
   "01111001100011" when "11101100",
   "01111001111001" when "11101101",
   "01111010001111" when "11101110",
   "01111010100101" when "11101111",
   "01111010111010" when "11110000",
   "01111011010000" when "11110001",
   "01111011100101" when "11110010",
   "01111011111011" when "11110011",
   "01111100010000" when "11110100",
   "01111100100101" when "11110101",
   "01111100111011" when "11110110",
   "01111101010000" when "11110111",
   "01111101100101" when "11111000",
   "01111101111010" when "11111001",
   "01111110001111" when "11111010",
   "01111110100011" when "11111011",
   "01111110111000" when "11111100",
   "01111111001101" when "11111101",
   "01111111100001" when "11111110",
   "01111111110110" when "11111111",
   "--------------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                        GenericTable_9_6_F400_uid33
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity GenericTable_9_6_F400_uid33 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(8 downto 0);
          Y : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of GenericTable_9_6_F400_uid33 is
signal TableOut :  std_logic_vector(5 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
  with X select TableOut <= 
   "101100" when "000000000",
   "101101" when "000000001",
   "101101" when "000000010",
   "101110" when "000000011",
   "101111" when "000000100",
   "101111" when "000000101",
   "110000" when "000000110",
   "110000" when "000000111",
   "110001" when "000001000",
   "110010" when "000001001",
   "110010" when "000001010",
   "110011" when "000001011",
   "110100" when "000001100",
   "110100" when "000001101",
   "110101" when "000001110",
   "110110" when "000001111",
   "110110" when "000010000",
   "110111" when "000010001",
   "110111" when "000010010",
   "111000" when "000010011",
   "111001" when "000010100",
   "111001" when "000010101",
   "111010" when "000010110",
   "111011" when "000010111",
   "111011" when "000011000",
   "111100" when "000011001",
   "111101" when "000011010",
   "111101" when "000011011",
   "111110" when "000011100",
   "111110" when "000011101",
   "111111" when "000011110",
   "111111" when "000011111",
   "101100" when "000100000",
   "101101" when "000100001",
   "101101" when "000100010",
   "101110" when "000100011",
   "101111" when "000100100",
   "101111" when "000100101",
   "110000" when "000100110",
   "110001" when "000100111",
   "110001" when "000101000",
   "110010" when "000101001",
   "110010" when "000101010",
   "110011" when "000101011",
   "110100" when "000101100",
   "110100" when "000101101",
   "110101" when "000101110",
   "110110" when "000101111",
   "110110" when "000110000",
   "110111" when "000110001",
   "110111" when "000110010",
   "111000" when "000110011",
   "111001" when "000110100",
   "111001" when "000110101",
   "111010" when "000110110",
   "111011" when "000110111",
   "111011" when "000111000",
   "111100" when "000111001",
   "111101" when "000111010",
   "111101" when "000111011",
   "111110" when "000111100",
   "111110" when "000111101",
   "111111" when "000111110",
   "111111" when "000111111",
   "101100" when "001000000",
   "101101" when "001000001",
   "101110" when "001000010",
   "101110" when "001000011",
   "101111" when "001000100",
   "110000" when "001000101",
   "110000" when "001000110",
   "110001" when "001000111",
   "110001" when "001001000",
   "110010" when "001001001",
   "110011" when "001001010",
   "110011" when "001001011",
   "110100" when "001001100",
   "110101" when "001001101",
   "110101" when "001001110",
   "110110" when "001001111",
   "110110" when "001010000",
   "110111" when "001010001",
   "111000" when "001010010",
   "111000" when "001010011",
   "111001" when "001010100",
   "111001" when "001010101",
   "111010" when "001010110",
   "111011" when "001010111",
   "111011" when "001011000",
   "111100" when "001011001",
   "111101" when "001011010",
   "111101" when "001011011",
   "111110" when "001011100",
   "111110" when "001011101",
   "111111" when "001011110",
   "111111" when "001011111",
   "101101" when "001100000",
   "101101" when "001100001",
   "101110" when "001100010",
   "101111" when "001100011",
   "101111" when "001100100",
   "110000" when "001100101",
   "110001" when "001100110",
   "110001" when "001100111",
   "110010" when "001101000",
   "110010" when "001101001",
   "110011" when "001101010",
   "110100" when "001101011",
   "110100" when "001101100",
   "110101" when "001101101",
   "110101" when "001101110",
   "110110" when "001101111",
   "110111" when "001110000",
   "110111" when "001110001",
   "111000" when "001110010",
   "111000" when "001110011",
   "111001" when "001110100",
   "111010" when "001110101",
   "111010" when "001110110",
   "111011" when "001110111",
   "111011" when "001111000",
   "111100" when "001111001",
   "111101" when "001111010",
   "111101" when "001111011",
   "111110" when "001111100",
   "111110" when "001111101",
   "111111" when "001111110",
   "111111" when "001111111",
   "101101" when "010000000",
   "101110" when "010000001",
   "101111" when "010000010",
   "101111" when "010000011",
   "110000" when "010000100",
   "110000" when "010000101",
   "110001" when "010000110",
   "110010" when "010000111",
   "110010" when "010001000",
   "110011" when "010001001",
   "110011" when "010001010",
   "110100" when "010001011",
   "110100" when "010001100",
   "110101" when "010001101",
   "110110" when "010001110",
   "110110" when "010001111",
   "110111" when "010010000",
   "110111" when "010010001",
   "111000" when "010010010",
   "111001" when "010010011",
   "111001" when "010010100",
   "111010" when "010010101",
   "111010" when "010010110",
   "111011" when "010010111",
   "111100" when "010011000",
   "111100" when "010011001",
   "111101" when "010011010",
   "111101" when "010011011",
   "111110" when "010011100",
   "111111" when "010011101",
   "111111" when "010011110",
   "111111" when "010011111",
   "101110" when "010100000",
   "101111" when "010100001",
   "101111" when "010100010",
   "110000" when "010100011",
   "110000" when "010100100",
   "110001" when "010100101",
   "110001" when "010100110",
   "110010" when "010100111",
   "110011" when "010101000",
   "110011" when "010101001",
   "110100" when "010101010",
   "110100" when "010101011",
   "110101" when "010101100",
   "110101" when "010101101",
   "110110" when "010101110",
   "110111" when "010101111",
   "110111" when "010110000",
   "111000" when "010110001",
   "111000" when "010110010",
   "111001" when "010110011",
   "111001" when "010110100",
   "111010" when "010110101",
   "111011" when "010110110",
   "111011" when "010110111",
   "111100" when "010111000",
   "111100" when "010111001",
   "111101" when "010111010",
   "111101" when "010111011",
   "111110" when "010111100",
   "111111" when "010111101",
   "111111" when "010111110",
   "111111" when "010111111",
   "101111" when "011000000",
   "101111" when "011000001",
   "110000" when "011000010",
   "110000" when "011000011",
   "110001" when "011000100",
   "110010" when "011000101",
   "110010" when "011000110",
   "110011" when "011000111",
   "110011" when "011001000",
   "110100" when "011001001",
   "110100" when "011001010",
   "110101" when "011001011",
   "110101" when "011001100",
   "110110" when "011001101",
   "110110" when "011001110",
   "110111" when "011001111",
   "111000" when "011010000",
   "111000" when "011010001",
   "111001" when "011010010",
   "111001" when "011010011",
   "111010" when "011010100",
   "111010" when "011010101",
   "111011" when "011010110",
   "111011" when "011010111",
   "111100" when "011011000",
   "111100" when "011011001",
   "111101" when "011011010",
   "111110" when "011011011",
   "111110" when "011011100",
   "111111" when "011011101",
   "111111" when "011011110",
   "111111" when "011011111",
   "110000" when "011100000",
   "110000" when "011100001",
   "110001" when "011100010",
   "110001" when "011100011",
   "110010" when "011100100",
   "110010" when "011100101",
   "110011" when "011100110",
   "110011" when "011100111",
   "110100" when "011101000",
   "110100" when "011101001",
   "110101" when "011101010",
   "110101" when "011101011",
   "110110" when "011101100",
   "110110" when "011101101",
   "110111" when "011101110",
   "110111" when "011101111",
   "111000" when "011110000",
   "111000" when "011110001",
   "111001" when "011110010",
   "111001" when "011110011",
   "111010" when "011110100",
   "111011" when "011110101",
   "111011" when "011110110",
   "111100" when "011110111",
   "111100" when "011111000",
   "111101" when "011111001",
   "111101" when "011111010",
   "111110" when "011111011",
   "111110" when "011111100",
   "111111" when "011111101",
   "111111" when "011111110",
   "111111" when "011111111",
   "110000" when "100000000",
   "110001" when "100000001",
   "110001" when "100000010",
   "110010" when "100000011",
   "110010" when "100000100",
   "110011" when "100000101",
   "110011" when "100000110",
   "110100" when "100000111",
   "110100" when "100001000",
   "110101" when "100001001",
   "110101" when "100001010",
   "110110" when "100001011",
   "110110" when "100001100",
   "110111" when "100001101",
   "110111" when "100001110",
   "111000" when "100001111",
   "111000" when "100010000",
   "111001" when "100010001",
   "111001" when "100010010",
   "111010" when "100010011",
   "111010" when "100010100",
   "111011" when "100010101",
   "111011" when "100010110",
   "111100" when "100010111",
   "111100" when "100011000",
   "111101" when "100011001",
   "111101" when "100011010",
   "111110" when "100011011",
   "111110" when "100011100",
   "111111" when "100011101",
   "111111" when "100011110",
   "111111" when "100011111",
   "110001" when "100100000",
   "110010" when "100100001",
   "110010" when "100100010",
   "110011" when "100100011",
   "110011" when "100100100",
   "110100" when "100100101",
   "110100" when "100100110",
   "110100" when "100100111",
   "110101" when "100101000",
   "110101" when "100101001",
   "110110" when "100101010",
   "110110" when "100101011",
   "110111" when "100101100",
   "110111" when "100101101",
   "111000" when "100101110",
   "111000" when "100101111",
   "111001" when "100110000",
   "111001" when "100110001",
   "111010" when "100110010",
   "111010" when "100110011",
   "111011" when "100110100",
   "111011" when "100110101",
   "111100" when "100110110",
   "111100" when "100110111",
   "111100" when "100111000",
   "111101" when "100111001",
   "111101" when "100111010",
   "111110" when "100111011",
   "111110" when "100111100",
   "111111" when "100111101",
   "111111" when "100111110",
   "111111" when "100111111",
   "110010" when "101000000",
   "110010" when "101000001",
   "110011" when "101000010",
   "110011" when "101000011",
   "110100" when "101000100",
   "110100" when "101000101",
   "110101" when "101000110",
   "110101" when "101000111",
   "110110" when "101001000",
   "110110" when "101001001",
   "110110" when "101001010",
   "110111" when "101001011",
   "110111" when "101001100",
   "111000" when "101001101",
   "111000" when "101001110",
   "111001" when "101001111",
   "111001" when "101010000",
   "111010" when "101010001",
   "111010" when "101010010",
   "111010" when "101010011",
   "111011" when "101010100",
   "111011" when "101010101",
   "111100" when "101010110",
   "111100" when "101010111",
   "111101" when "101011000",
   "111101" when "101011001",
   "111110" when "101011010",
   "111110" when "101011011",
   "111110" when "101011100",
   "111111" when "101011101",
   "111111" when "101011110",
   "111111" when "101011111",
   "110011" when "101100000",
   "110011" when "101100001",
   "110100" when "101100010",
   "110100" when "101100011",
   "110100" when "101100100",
   "110101" when "101100101",
   "110101" when "101100110",
   "110110" when "101100111",
   "110110" when "101101000",
   "110111" when "101101001",
   "110111" when "101101010",
   "110111" when "101101011",
   "111000" when "101101100",
   "111000" when "101101101",
   "111001" when "101101110",
   "111001" when "101101111",
   "111001" when "101110000",
   "111010" when "101110001",
   "111010" when "101110010",
   "111011" when "101110011",
   "111011" when "101110100",
   "111100" when "101110101",
   "111100" when "101110110",
   "111100" when "101110111",
   "111101" when "101111000",
   "111101" when "101111001",
   "111110" when "101111010",
   "111110" when "101111011",
   "111111" when "101111100",
   "111111" when "101111101",
   "111111" when "101111110",
   "111111" when "101111111",
   "110100" when "110000000",
   "110100" when "110000001",
   "110100" when "110000010",
   "110101" when "110000011",
   "110101" when "110000100",
   "110110" when "110000101",
   "110110" when "110000110",
   "110110" when "110000111",
   "110111" when "110001000",
   "110111" when "110001001",
   "111000" when "110001010",
   "111000" when "110001011",
   "111000" when "110001100",
   "111001" when "110001101",
   "111001" when "110001110",
   "111001" when "110001111",
   "111010" when "110010000",
   "111010" when "110010001",
   "111011" when "110010010",
   "111011" when "110010011",
   "111011" when "110010100",
   "111100" when "110010101",
   "111100" when "110010110",
   "111101" when "110010111",
   "111101" when "110011000",
   "111101" when "110011001",
   "111110" when "110011010",
   "111110" when "110011011",
   "111111" when "110011100",
   "111111" when "110011101",
   "111111" when "110011110",
   "111111" when "110011111",
   "110100" when "110100000",
   "110101" when "110100001",
   "110101" when "110100010",
   "110101" when "110100011",
   "110110" when "110100100",
   "110110" when "110100101",
   "110111" when "110100110",
   "110111" when "110100111",
   "110111" when "110101000",
   "111000" when "110101001",
   "111000" when "110101010",
   "111000" when "110101011",
   "111001" when "110101100",
   "111001" when "110101101",
   "111001" when "110101110",
   "111010" when "110101111",
   "111010" when "110110000",
   "111011" when "110110001",
   "111011" when "110110010",
   "111011" when "110110011",
   "111100" when "110110100",
   "111100" when "110110101",
   "111100" when "110110110",
   "111101" when "110110111",
   "111101" when "110111000",
   "111110" when "110111001",
   "111110" when "110111010",
   "111110" when "110111011",
   "111111" when "110111100",
   "111111" when "110111101",
   "111111" when "110111110",
   "111111" when "110111111",
   "110101" when "111000000",
   "110101" when "111000001",
   "110110" when "111000010",
   "110110" when "111000011",
   "110110" when "111000100",
   "110111" when "111000101",
   "110111" when "111000110",
   "110111" when "111000111",
   "111000" when "111001000",
   "111000" when "111001001",
   "111000" when "111001010",
   "111001" when "111001011",
   "111001" when "111001100",
   "111010" when "111001101",
   "111010" when "111001110",
   "111010" when "111001111",
   "111011" when "111010000",
   "111011" when "111010001",
   "111011" when "111010010",
   "111100" when "111010011",
   "111100" when "111010100",
   "111100" when "111010101",
   "111101" when "111010110",
   "111101" when "111010111",
   "111101" when "111011000",
   "111110" when "111011001",
   "111110" when "111011010",
   "111110" when "111011011",
   "111111" when "111011100",
   "111111" when "111011101",
   "111111" when "111011110",
   "111111" when "111011111",
   "110110" when "111100000",
   "110110" when "111100001",
   "110110" when "111100010",
   "110111" when "111100011",
   "110111" when "111100100",
   "110111" when "111100101",
   "111000" when "111100110",
   "111000" when "111100111",
   "111000" when "111101000",
   "111001" when "111101001",
   "111001" when "111101010",
   "111001" when "111101011",
   "111010" when "111101100",
   "111010" when "111101101",
   "111010" when "111101110",
   "111011" when "111101111",
   "111011" when "111110000",
   "111011" when "111110001",
   "111100" when "111110010",
   "111100" when "111110011",
   "111100" when "111110100",
   "111101" when "111110101",
   "111101" when "111110110",
   "111101" when "111110111",
   "111110" when "111111000",
   "111110" when "111111001",
   "111110" when "111111010",
   "111111" when "111111011",
   "111111" when "111111100",
   "111111" when "111111101",
   "111111" when "111111110",
   "111111" when "111111111",
   "------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                                 atan_uid36
--         (BipartiteTable_f_atan_x_pi_in_M14_out_M2_M13_F400_uid27)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Matei Istoan (2014)
--------------------------------------------------------------------------------
-- Pipeline depth: 0 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity atan_uid36 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(13 downto 0);
          Y : out  std_logic_vector(11 downto 0)   );
end entity;

architecture arch of atan_uid36 is
   component GenericTable_8_14_F400_uid29 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(7 downto 0);
             Y : out  std_logic_vector(13 downto 0)   );
   end component;

   component GenericTable_9_6_F400_uid33 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(8 downto 0);
             Y : out  std_logic_vector(5 downto 0)   );
   end component;

signal X0 :  std_logic_vector(3 downto 0);
signal X1 :  std_logic_vector(3 downto 0);
signal X2 :  std_logic_vector(5 downto 0);
signal X2_msb :  std_logic;
signal X2_short :  std_logic_vector(4 downto 0);
signal X2_short_inv :  std_logic_vector(4 downto 0);
signal tableTIVaddr :  std_logic_vector(7 downto 0);
signal tableTOaddr :  std_logic_vector(8 downto 0);
signal tableTIVout :  std_logic_vector(13 downto 0);
signal tableTOout :  std_logic_vector(5 downto 0);
signal tableTOout_inv :  std_logic_vector(5 downto 0);
signal tableTIV_fxp :  signed(-2+15 downto 0);
signal tableTO_fxp :  signed(-10+15 downto 0);
signal tableTO_fxp_sgnExt :  signed(-2+15 downto 0);
signal Y_int :  signed(-2+15 downto 0);
signal Y_int_short :  signed(-2+14 downto 0);
signal Y_rnd :  signed(-2+14 downto 0);
attribute rom_extract: string;
attribute rom_style: string;
attribute rom_extract of GenericTable_8_14_F400_uid29: component is "yes";
attribute rom_extract of GenericTable_9_6_F400_uid33: component is "yes";
attribute rom_style of GenericTable_8_14_F400_uid29: component is "block";
attribute rom_style of GenericTable_9_6_F400_uid33: component is "block";
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
         end if;
      end process;
   X0 <= X(13 downto 10);
   X1 <= X(9 downto 6);
   X2 <= X(5 downto 0);

   X2_msb <= X2(5);
   X2_short <= X2(4 downto 0);
   X2_short_inv <= X2_short xor (4 downto 0 => X2_msb);

   tableTIVaddr <= X0 & X1;
   tableTOaddr <= X0 & X2_short_inv;

   TIVtable: GenericTable_8_14_F400_uid29  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => tableTIVaddr,
                 Y => tableTIVout);

   TOtable: GenericTable_9_6_F400_uid33  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => tableTOaddr,
                 Y => tableTOout);

   tableTOout_inv <= tableTOout xor (5 downto 0 => X2_msb);

   tableTIV_fxp <= signed(tableTIVout);
   tableTO_fxp <= signed(tableTOout_inv);
   tableTO_fxp_sgnExt <= (7 downto 0 => tableTO_fxp(5)) & tableTO_fxp(5 downto 0); -- fix resize from (-10, -15) to (-2, -15)

   Y_int <= tableTIV_fxp + tableTO_fxp_sgnExt;
   Y_int_short <= Y_int(13 downto 1); -- fix resize from (-2, -15) to (-2, -14)
   Y_rnd <= Y_int_short + ("000000000000" & '1');
   Y <= std_logic_vector(Y_rnd(12 downto 1));
end architecture;

--------------------------------------------------------------------------------
--                  FixAtan2ByRecipMultAtan_14_14_F400_uid2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Matei Istoan, Florent de Dinechin (2012-...)
--------------------------------------------------------------------------------
-- Pipeline depth: 4 cycles

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FixAtan2ByRecipMultAtan_14_14_F400_uid2 is
   port ( clk, rst : in std_logic;
          X : in  std_logic_vector(13 downto 0);
          Y : in  std_logic_vector(13 downto 0);
          A : out  std_logic_vector(13 downto 0)   );
end entity;

architecture arch of FixAtan2ByRecipMultAtan_14_14_F400_uid2 is
   component LZOC_12_F400_uid4 is
      port ( clk, rst : in std_logic;
             I : in  std_logic_vector(11 downto 0);
             OZB : in  std_logic;
             O : out  std_logic_vector(3 downto 0)   );
   end component;

   component LeftShifter_13_by_max_12_F400_uid8 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(12 downto 0);
             S : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(24 downto 0)   );
   end component;

   component reciprocal_uid23 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(11 downto 0);
             Y : out  std_logic_vector(15 downto 0)   );
   end component;

   component atan_uid36 is
      port ( clk, rst : in std_logic;
             X : in  std_logic_vector(13 downto 0);
             Y : out  std_logic_vector(11 downto 0)   );
   end component;

signal sgnX :  std_logic;
signal sgnY :  std_logic;
signal Xsat :  std_logic_vector(13 downto 0);
signal Ysat :  std_logic_vector(13 downto 0);
signal pX :  std_logic_vector(13 downto 0);
signal pY :  std_logic_vector(13 downto 0);
signal mX :  std_logic_vector(13 downto 0);
signal mY :  std_logic_vector(13 downto 0);
signal XmY :  std_logic_vector(14 downto 0);
signal XpY :  std_logic_vector(14 downto 0);
signal XltY :  std_logic;
signal mYltX :  std_logic;
signal quadrant, quadrant_d1, quadrant_d2, quadrant_d3, quadrant_d4 :  std_logic_vector(1 downto 0);
signal XR, XR_d1, XR_d2 :  std_logic_vector(12 downto 0);
signal YR, YR_d1, YR_d2 :  std_logic_vector(12 downto 0);
signal finalAdd, finalAdd_d1, finalAdd_d2, finalAdd_d3, finalAdd_d4 :  std_logic;
signal XorY :  std_logic_vector(11 downto 0);
signal S :  std_logic_vector(3 downto 0);
signal XRSfull :  std_logic_vector(24 downto 0);
signal XRS, XRS_d1 :  std_logic_vector(12 downto 0);
signal YRSfull :  std_logic_vector(24 downto 0);
signal YRS, YRS_d1 :  std_logic_vector(12 downto 0);
signal XRm1 :  std_logic_vector(11 downto 0);
signal R0 :  std_logic_vector(15 downto 0);
signal R, R_d1 :  unsigned(0+14 downto 0);
signal YRU, YRU_d1 :  unsigned(-1+13 downto 0);
signal P :  unsigned(0+27 downto 0);
signal PtruncU :  unsigned(-1+14 downto 0);
signal P_slv :  std_logic_vector(13 downto 0);
signal atanTableOut :  std_logic_vector(11 downto 0);
signal finalZ :  std_logic_vector(13 downto 0);
signal qangle :  std_logic_vector(13 downto 0);
begin
   process(clk)
      begin
         if clk'event and clk = '1' then
            quadrant_d1 <=  quadrant;
            quadrant_d2 <=  quadrant_d1;
            quadrant_d3 <=  quadrant_d2;
            quadrant_d4 <=  quadrant_d3;
            XR_d1 <=  XR;
            XR_d2 <=  XR_d1;
            YR_d1 <=  YR;
            YR_d2 <=  YR_d1;
            finalAdd_d1 <=  finalAdd;
            finalAdd_d2 <=  finalAdd_d1;
            finalAdd_d3 <=  finalAdd_d2;
            finalAdd_d4 <=  finalAdd_d3;
            XRS_d1 <=  XRS;
            YRS_d1 <=  YRS;
            R_d1 <=  R;
            YRU_d1 <=  YRU;
         end if;
      end process;
   sgnX <= X(13);
   sgnY <= Y(13);
   -- First saturate x and y in case they touch -1
   Xsat <= "10000000000001" when X="10000000000000" else X ;
   Ysat <= "10000000000001" when Y="10000000000000" else Y ;
   pX <= Xsat;
   pY <= Ysat;
   mX <= ("00000000000000" - Xsat);
   mY <= ("00000000000000" - Ysat);
   XmY <= (sgnX & Xsat)-(sgnY & Ysat);
   XpY <= (sgnX & Xsat)+(sgnY & Ysat);
   XltY <= XmY(14);
   mYltX <= not XpY(14);
   -- quadrant will also be the angle to add at the end
   quadrant <= 
      "00"  when (not sgnX and not XltY and     mYltX)='1' else
      "01"  when (not sgnY and     XltY and     mYltX)='1' else
      "10"  when (    sgnX and     XltY and not mYltX)='1' else
      "11";
   XR <= 
      pX(12 downto 0) when quadrant="00"   else 
      pY(12 downto 0) when quadrant="01"   else 
      mX(12 downto 0) when quadrant="10"   else 
      mY(12 downto 0);
   YR <= 
      pY(12 downto 0) when quadrant="00" and sgnY='0'  else 
      mY(12 downto 0) when quadrant="00" and sgnY='1'  else 
      pX(12 downto 0) when quadrant="01" and sgnX='0'  else 
      mX(12 downto 0) when quadrant="01" and sgnX='1'  else 
      pY(12 downto 0) when quadrant="10" and sgnY='0'  else 
      mY(12 downto 0) when quadrant="10" and sgnY='1'  else 
      pX(12 downto 0) when quadrant="11" and sgnX='0'  else 
      mX(12 downto 0) ;
   finalAdd <= 
      '1' when (quadrant="00" and sgnY='0') or(quadrant="01" and sgnX='1') or (quadrant="10" and sgnY='1') or (quadrant="11" and sgnX='0')
       else '0';  -- this information is sent to the end of the pipeline, better compute it here as one bit
   XorY <= XR(12 downto 1) or YR(12 downto 1);
   lzc: LZOC_12_F400_uid4  -- pipelineDepth=2 maxInDelay=2.05144e-09
      port map ( clk  => clk,
                 rst  => rst,
                 I => XorY,
                 O => S,
                 OZB => '0');
   ----------------Synchro barrier, entering cycle 2----------------
   Xshift: LeftShifter_13_by_max_12_F400_uid8  -- pipelineDepth=1 maxInDelay=1.07033e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => XRSfull,
                 S => S,
                 X => XR_d2);
   XRS <=  XRSfull (12 downto 0);
   Yshift: LeftShifter_13_by_max_12_F400_uid8  -- pipelineDepth=1 maxInDelay=1.07033e-09
      port map ( clk  => clk,
                 rst  => rst,
                 R => YRSfull,
                 S => S,
                 X => YR_d2);
   YRS <=  YRSfull (12 downto 0);
   ----------------Synchro barrier, entering cycle 3----------------
   XRm1 <= XRS_d1(11 downto 0); -- removing the MSB which is constantly 1
   recipTable: reciprocal_uid23  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => XRm1,
                 Y => R0);
   R <= unsigned(R0(14 downto 0)); -- removing the sign  bit
   YRU <= unsigned(YRS_d1);
   ----------------Synchro barrier, entering cycle 4----------------
   P <= R_d1*YRU_d1;
   PtruncU <= P(26 downto 13); -- fix resize from (0, -27) to (-1, -14)
   P_slv <=  std_logic_vector(PtruncU);
   atanTable: atan_uid36  -- pipelineDepth=0 maxInDelay=0
      port map ( clk  => clk,
                 rst  => rst,
                 X => P_slv,
                 Y => atanTableOut);
   finalZ <= "00" & atanTableOut;
   qangle <= (quadrant_d4 & "000000000000");
   A <=            qangle + finalZ  when finalAdd_d4='1'
      else qangle - finalZ;
end architecture;

